module mem_0_ext(
  input  [33:0] R0_addr,
  input         R0_clk,
  output [63:0] R0_data,
  input         R0_en,
  input  [33:0] W0_addr,
  input         W0_clk,
  input  [63:0] W0_data,
  input         W0_en,
  input  [7:0]  W0_mask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire [25:0] mem_0_0_R0_addr;
  wire  mem_0_0_R0_clk;
  wire [7:0] mem_0_0_R0_data;
  wire  mem_0_0_R0_en;
  wire [25:0] mem_0_0_W0_addr;
  wire  mem_0_0_W0_clk;
  wire [7:0] mem_0_0_W0_data;
  wire  mem_0_0_W0_en;
  wire  mem_0_0_W0_mask;
  wire [25:0] mem_0_1_R0_addr;
  wire  mem_0_1_R0_clk;
  wire [7:0] mem_0_1_R0_data;
  wire  mem_0_1_R0_en;
  wire [25:0] mem_0_1_W0_addr;
  wire  mem_0_1_W0_clk;
  wire [7:0] mem_0_1_W0_data;
  wire  mem_0_1_W0_en;
  wire  mem_0_1_W0_mask;
  wire [25:0] mem_0_2_R0_addr;
  wire  mem_0_2_R0_clk;
  wire [7:0] mem_0_2_R0_data;
  wire  mem_0_2_R0_en;
  wire [25:0] mem_0_2_W0_addr;
  wire  mem_0_2_W0_clk;
  wire [7:0] mem_0_2_W0_data;
  wire  mem_0_2_W0_en;
  wire  mem_0_2_W0_mask;
  wire [25:0] mem_0_3_R0_addr;
  wire  mem_0_3_R0_clk;
  wire [7:0] mem_0_3_R0_data;
  wire  mem_0_3_R0_en;
  wire [25:0] mem_0_3_W0_addr;
  wire  mem_0_3_W0_clk;
  wire [7:0] mem_0_3_W0_data;
  wire  mem_0_3_W0_en;
  wire  mem_0_3_W0_mask;
  wire [25:0] mem_0_4_R0_addr;
  wire  mem_0_4_R0_clk;
  wire [7:0] mem_0_4_R0_data;
  wire  mem_0_4_R0_en;
  wire [25:0] mem_0_4_W0_addr;
  wire  mem_0_4_W0_clk;
  wire [7:0] mem_0_4_W0_data;
  wire  mem_0_4_W0_en;
  wire  mem_0_4_W0_mask;
  wire [25:0] mem_0_5_R0_addr;
  wire  mem_0_5_R0_clk;
  wire [7:0] mem_0_5_R0_data;
  wire  mem_0_5_R0_en;
  wire [25:0] mem_0_5_W0_addr;
  wire  mem_0_5_W0_clk;
  wire [7:0] mem_0_5_W0_data;
  wire  mem_0_5_W0_en;
  wire  mem_0_5_W0_mask;
  wire [25:0] mem_0_6_R0_addr;
  wire  mem_0_6_R0_clk;
  wire [7:0] mem_0_6_R0_data;
  wire  mem_0_6_R0_en;
  wire [25:0] mem_0_6_W0_addr;
  wire  mem_0_6_W0_clk;
  wire [7:0] mem_0_6_W0_data;
  wire  mem_0_6_W0_en;
  wire  mem_0_6_W0_mask;
  wire [25:0] mem_0_7_R0_addr;
  wire  mem_0_7_R0_clk;
  wire [7:0] mem_0_7_R0_data;
  wire  mem_0_7_R0_en;
  wire [25:0] mem_0_7_W0_addr;
  wire  mem_0_7_W0_clk;
  wire [7:0] mem_0_7_W0_data;
  wire  mem_0_7_W0_en;
  wire  mem_0_7_W0_mask;
  wire [25:0] mem_1_0_R0_addr;
  wire  mem_1_0_R0_clk;
  wire [7:0] mem_1_0_R0_data;
  wire  mem_1_0_R0_en;
  wire [25:0] mem_1_0_W0_addr;
  wire  mem_1_0_W0_clk;
  wire [7:0] mem_1_0_W0_data;
  wire  mem_1_0_W0_en;
  wire  mem_1_0_W0_mask;
  wire [25:0] mem_1_1_R0_addr;
  wire  mem_1_1_R0_clk;
  wire [7:0] mem_1_1_R0_data;
  wire  mem_1_1_R0_en;
  wire [25:0] mem_1_1_W0_addr;
  wire  mem_1_1_W0_clk;
  wire [7:0] mem_1_1_W0_data;
  wire  mem_1_1_W0_en;
  wire  mem_1_1_W0_mask;
  wire [25:0] mem_1_2_R0_addr;
  wire  mem_1_2_R0_clk;
  wire [7:0] mem_1_2_R0_data;
  wire  mem_1_2_R0_en;
  wire [25:0] mem_1_2_W0_addr;
  wire  mem_1_2_W0_clk;
  wire [7:0] mem_1_2_W0_data;
  wire  mem_1_2_W0_en;
  wire  mem_1_2_W0_mask;
  wire [25:0] mem_1_3_R0_addr;
  wire  mem_1_3_R0_clk;
  wire [7:0] mem_1_3_R0_data;
  wire  mem_1_3_R0_en;
  wire [25:0] mem_1_3_W0_addr;
  wire  mem_1_3_W0_clk;
  wire [7:0] mem_1_3_W0_data;
  wire  mem_1_3_W0_en;
  wire  mem_1_3_W0_mask;
  wire [25:0] mem_1_4_R0_addr;
  wire  mem_1_4_R0_clk;
  wire [7:0] mem_1_4_R0_data;
  wire  mem_1_4_R0_en;
  wire [25:0] mem_1_4_W0_addr;
  wire  mem_1_4_W0_clk;
  wire [7:0] mem_1_4_W0_data;
  wire  mem_1_4_W0_en;
  wire  mem_1_4_W0_mask;
  wire [25:0] mem_1_5_R0_addr;
  wire  mem_1_5_R0_clk;
  wire [7:0] mem_1_5_R0_data;
  wire  mem_1_5_R0_en;
  wire [25:0] mem_1_5_W0_addr;
  wire  mem_1_5_W0_clk;
  wire [7:0] mem_1_5_W0_data;
  wire  mem_1_5_W0_en;
  wire  mem_1_5_W0_mask;
  wire [25:0] mem_1_6_R0_addr;
  wire  mem_1_6_R0_clk;
  wire [7:0] mem_1_6_R0_data;
  wire  mem_1_6_R0_en;
  wire [25:0] mem_1_6_W0_addr;
  wire  mem_1_6_W0_clk;
  wire [7:0] mem_1_6_W0_data;
  wire  mem_1_6_W0_en;
  wire  mem_1_6_W0_mask;
  wire [25:0] mem_1_7_R0_addr;
  wire  mem_1_7_R0_clk;
  wire [7:0] mem_1_7_R0_data;
  wire  mem_1_7_R0_en;
  wire [25:0] mem_1_7_W0_addr;
  wire  mem_1_7_W0_clk;
  wire [7:0] mem_1_7_W0_data;
  wire  mem_1_7_W0_en;
  wire  mem_1_7_W0_mask;
  wire [25:0] mem_2_0_R0_addr;
  wire  mem_2_0_R0_clk;
  wire [7:0] mem_2_0_R0_data;
  wire  mem_2_0_R0_en;
  wire [25:0] mem_2_0_W0_addr;
  wire  mem_2_0_W0_clk;
  wire [7:0] mem_2_0_W0_data;
  wire  mem_2_0_W0_en;
  wire  mem_2_0_W0_mask;
  wire [25:0] mem_2_1_R0_addr;
  wire  mem_2_1_R0_clk;
  wire [7:0] mem_2_1_R0_data;
  wire  mem_2_1_R0_en;
  wire [25:0] mem_2_1_W0_addr;
  wire  mem_2_1_W0_clk;
  wire [7:0] mem_2_1_W0_data;
  wire  mem_2_1_W0_en;
  wire  mem_2_1_W0_mask;
  wire [25:0] mem_2_2_R0_addr;
  wire  mem_2_2_R0_clk;
  wire [7:0] mem_2_2_R0_data;
  wire  mem_2_2_R0_en;
  wire [25:0] mem_2_2_W0_addr;
  wire  mem_2_2_W0_clk;
  wire [7:0] mem_2_2_W0_data;
  wire  mem_2_2_W0_en;
  wire  mem_2_2_W0_mask;
  wire [25:0] mem_2_3_R0_addr;
  wire  mem_2_3_R0_clk;
  wire [7:0] mem_2_3_R0_data;
  wire  mem_2_3_R0_en;
  wire [25:0] mem_2_3_W0_addr;
  wire  mem_2_3_W0_clk;
  wire [7:0] mem_2_3_W0_data;
  wire  mem_2_3_W0_en;
  wire  mem_2_3_W0_mask;
  wire [25:0] mem_2_4_R0_addr;
  wire  mem_2_4_R0_clk;
  wire [7:0] mem_2_4_R0_data;
  wire  mem_2_4_R0_en;
  wire [25:0] mem_2_4_W0_addr;
  wire  mem_2_4_W0_clk;
  wire [7:0] mem_2_4_W0_data;
  wire  mem_2_4_W0_en;
  wire  mem_2_4_W0_mask;
  wire [25:0] mem_2_5_R0_addr;
  wire  mem_2_5_R0_clk;
  wire [7:0] mem_2_5_R0_data;
  wire  mem_2_5_R0_en;
  wire [25:0] mem_2_5_W0_addr;
  wire  mem_2_5_W0_clk;
  wire [7:0] mem_2_5_W0_data;
  wire  mem_2_5_W0_en;
  wire  mem_2_5_W0_mask;
  wire [25:0] mem_2_6_R0_addr;
  wire  mem_2_6_R0_clk;
  wire [7:0] mem_2_6_R0_data;
  wire  mem_2_6_R0_en;
  wire [25:0] mem_2_6_W0_addr;
  wire  mem_2_6_W0_clk;
  wire [7:0] mem_2_6_W0_data;
  wire  mem_2_6_W0_en;
  wire  mem_2_6_W0_mask;
  wire [25:0] mem_2_7_R0_addr;
  wire  mem_2_7_R0_clk;
  wire [7:0] mem_2_7_R0_data;
  wire  mem_2_7_R0_en;
  wire [25:0] mem_2_7_W0_addr;
  wire  mem_2_7_W0_clk;
  wire [7:0] mem_2_7_W0_data;
  wire  mem_2_7_W0_en;
  wire  mem_2_7_W0_mask;
  wire [25:0] mem_3_0_R0_addr;
  wire  mem_3_0_R0_clk;
  wire [7:0] mem_3_0_R0_data;
  wire  mem_3_0_R0_en;
  wire [25:0] mem_3_0_W0_addr;
  wire  mem_3_0_W0_clk;
  wire [7:0] mem_3_0_W0_data;
  wire  mem_3_0_W0_en;
  wire  mem_3_0_W0_mask;
  wire [25:0] mem_3_1_R0_addr;
  wire  mem_3_1_R0_clk;
  wire [7:0] mem_3_1_R0_data;
  wire  mem_3_1_R0_en;
  wire [25:0] mem_3_1_W0_addr;
  wire  mem_3_1_W0_clk;
  wire [7:0] mem_3_1_W0_data;
  wire  mem_3_1_W0_en;
  wire  mem_3_1_W0_mask;
  wire [25:0] mem_3_2_R0_addr;
  wire  mem_3_2_R0_clk;
  wire [7:0] mem_3_2_R0_data;
  wire  mem_3_2_R0_en;
  wire [25:0] mem_3_2_W0_addr;
  wire  mem_3_2_W0_clk;
  wire [7:0] mem_3_2_W0_data;
  wire  mem_3_2_W0_en;
  wire  mem_3_2_W0_mask;
  wire [25:0] mem_3_3_R0_addr;
  wire  mem_3_3_R0_clk;
  wire [7:0] mem_3_3_R0_data;
  wire  mem_3_3_R0_en;
  wire [25:0] mem_3_3_W0_addr;
  wire  mem_3_3_W0_clk;
  wire [7:0] mem_3_3_W0_data;
  wire  mem_3_3_W0_en;
  wire  mem_3_3_W0_mask;
  wire [25:0] mem_3_4_R0_addr;
  wire  mem_3_4_R0_clk;
  wire [7:0] mem_3_4_R0_data;
  wire  mem_3_4_R0_en;
  wire [25:0] mem_3_4_W0_addr;
  wire  mem_3_4_W0_clk;
  wire [7:0] mem_3_4_W0_data;
  wire  mem_3_4_W0_en;
  wire  mem_3_4_W0_mask;
  wire [25:0] mem_3_5_R0_addr;
  wire  mem_3_5_R0_clk;
  wire [7:0] mem_3_5_R0_data;
  wire  mem_3_5_R0_en;
  wire [25:0] mem_3_5_W0_addr;
  wire  mem_3_5_W0_clk;
  wire [7:0] mem_3_5_W0_data;
  wire  mem_3_5_W0_en;
  wire  mem_3_5_W0_mask;
  wire [25:0] mem_3_6_R0_addr;
  wire  mem_3_6_R0_clk;
  wire [7:0] mem_3_6_R0_data;
  wire  mem_3_6_R0_en;
  wire [25:0] mem_3_6_W0_addr;
  wire  mem_3_6_W0_clk;
  wire [7:0] mem_3_6_W0_data;
  wire  mem_3_6_W0_en;
  wire  mem_3_6_W0_mask;
  wire [25:0] mem_3_7_R0_addr;
  wire  mem_3_7_R0_clk;
  wire [7:0] mem_3_7_R0_data;
  wire  mem_3_7_R0_en;
  wire [25:0] mem_3_7_W0_addr;
  wire  mem_3_7_W0_clk;
  wire [7:0] mem_3_7_W0_data;
  wire  mem_3_7_W0_en;
  wire  mem_3_7_W0_mask;
  wire [25:0] mem_4_0_R0_addr;
  wire  mem_4_0_R0_clk;
  wire [7:0] mem_4_0_R0_data;
  wire  mem_4_0_R0_en;
  wire [25:0] mem_4_0_W0_addr;
  wire  mem_4_0_W0_clk;
  wire [7:0] mem_4_0_W0_data;
  wire  mem_4_0_W0_en;
  wire  mem_4_0_W0_mask;
  wire [25:0] mem_4_1_R0_addr;
  wire  mem_4_1_R0_clk;
  wire [7:0] mem_4_1_R0_data;
  wire  mem_4_1_R0_en;
  wire [25:0] mem_4_1_W0_addr;
  wire  mem_4_1_W0_clk;
  wire [7:0] mem_4_1_W0_data;
  wire  mem_4_1_W0_en;
  wire  mem_4_1_W0_mask;
  wire [25:0] mem_4_2_R0_addr;
  wire  mem_4_2_R0_clk;
  wire [7:0] mem_4_2_R0_data;
  wire  mem_4_2_R0_en;
  wire [25:0] mem_4_2_W0_addr;
  wire  mem_4_2_W0_clk;
  wire [7:0] mem_4_2_W0_data;
  wire  mem_4_2_W0_en;
  wire  mem_4_2_W0_mask;
  wire [25:0] mem_4_3_R0_addr;
  wire  mem_4_3_R0_clk;
  wire [7:0] mem_4_3_R0_data;
  wire  mem_4_3_R0_en;
  wire [25:0] mem_4_3_W0_addr;
  wire  mem_4_3_W0_clk;
  wire [7:0] mem_4_3_W0_data;
  wire  mem_4_3_W0_en;
  wire  mem_4_3_W0_mask;
  wire [25:0] mem_4_4_R0_addr;
  wire  mem_4_4_R0_clk;
  wire [7:0] mem_4_4_R0_data;
  wire  mem_4_4_R0_en;
  wire [25:0] mem_4_4_W0_addr;
  wire  mem_4_4_W0_clk;
  wire [7:0] mem_4_4_W0_data;
  wire  mem_4_4_W0_en;
  wire  mem_4_4_W0_mask;
  wire [25:0] mem_4_5_R0_addr;
  wire  mem_4_5_R0_clk;
  wire [7:0] mem_4_5_R0_data;
  wire  mem_4_5_R0_en;
  wire [25:0] mem_4_5_W0_addr;
  wire  mem_4_5_W0_clk;
  wire [7:0] mem_4_5_W0_data;
  wire  mem_4_5_W0_en;
  wire  mem_4_5_W0_mask;
  wire [25:0] mem_4_6_R0_addr;
  wire  mem_4_6_R0_clk;
  wire [7:0] mem_4_6_R0_data;
  wire  mem_4_6_R0_en;
  wire [25:0] mem_4_6_W0_addr;
  wire  mem_4_6_W0_clk;
  wire [7:0] mem_4_6_W0_data;
  wire  mem_4_6_W0_en;
  wire  mem_4_6_W0_mask;
  wire [25:0] mem_4_7_R0_addr;
  wire  mem_4_7_R0_clk;
  wire [7:0] mem_4_7_R0_data;
  wire  mem_4_7_R0_en;
  wire [25:0] mem_4_7_W0_addr;
  wire  mem_4_7_W0_clk;
  wire [7:0] mem_4_7_W0_data;
  wire  mem_4_7_W0_en;
  wire  mem_4_7_W0_mask;
  wire [25:0] mem_5_0_R0_addr;
  wire  mem_5_0_R0_clk;
  wire [7:0] mem_5_0_R0_data;
  wire  mem_5_0_R0_en;
  wire [25:0] mem_5_0_W0_addr;
  wire  mem_5_0_W0_clk;
  wire [7:0] mem_5_0_W0_data;
  wire  mem_5_0_W0_en;
  wire  mem_5_0_W0_mask;
  wire [25:0] mem_5_1_R0_addr;
  wire  mem_5_1_R0_clk;
  wire [7:0] mem_5_1_R0_data;
  wire  mem_5_1_R0_en;
  wire [25:0] mem_5_1_W0_addr;
  wire  mem_5_1_W0_clk;
  wire [7:0] mem_5_1_W0_data;
  wire  mem_5_1_W0_en;
  wire  mem_5_1_W0_mask;
  wire [25:0] mem_5_2_R0_addr;
  wire  mem_5_2_R0_clk;
  wire [7:0] mem_5_2_R0_data;
  wire  mem_5_2_R0_en;
  wire [25:0] mem_5_2_W0_addr;
  wire  mem_5_2_W0_clk;
  wire [7:0] mem_5_2_W0_data;
  wire  mem_5_2_W0_en;
  wire  mem_5_2_W0_mask;
  wire [25:0] mem_5_3_R0_addr;
  wire  mem_5_3_R0_clk;
  wire [7:0] mem_5_3_R0_data;
  wire  mem_5_3_R0_en;
  wire [25:0] mem_5_3_W0_addr;
  wire  mem_5_3_W0_clk;
  wire [7:0] mem_5_3_W0_data;
  wire  mem_5_3_W0_en;
  wire  mem_5_3_W0_mask;
  wire [25:0] mem_5_4_R0_addr;
  wire  mem_5_4_R0_clk;
  wire [7:0] mem_5_4_R0_data;
  wire  mem_5_4_R0_en;
  wire [25:0] mem_5_4_W0_addr;
  wire  mem_5_4_W0_clk;
  wire [7:0] mem_5_4_W0_data;
  wire  mem_5_4_W0_en;
  wire  mem_5_4_W0_mask;
  wire [25:0] mem_5_5_R0_addr;
  wire  mem_5_5_R0_clk;
  wire [7:0] mem_5_5_R0_data;
  wire  mem_5_5_R0_en;
  wire [25:0] mem_5_5_W0_addr;
  wire  mem_5_5_W0_clk;
  wire [7:0] mem_5_5_W0_data;
  wire  mem_5_5_W0_en;
  wire  mem_5_5_W0_mask;
  wire [25:0] mem_5_6_R0_addr;
  wire  mem_5_6_R0_clk;
  wire [7:0] mem_5_6_R0_data;
  wire  mem_5_6_R0_en;
  wire [25:0] mem_5_6_W0_addr;
  wire  mem_5_6_W0_clk;
  wire [7:0] mem_5_6_W0_data;
  wire  mem_5_6_W0_en;
  wire  mem_5_6_W0_mask;
  wire [25:0] mem_5_7_R0_addr;
  wire  mem_5_7_R0_clk;
  wire [7:0] mem_5_7_R0_data;
  wire  mem_5_7_R0_en;
  wire [25:0] mem_5_7_W0_addr;
  wire  mem_5_7_W0_clk;
  wire [7:0] mem_5_7_W0_data;
  wire  mem_5_7_W0_en;
  wire  mem_5_7_W0_mask;
  wire [25:0] mem_6_0_R0_addr;
  wire  mem_6_0_R0_clk;
  wire [7:0] mem_6_0_R0_data;
  wire  mem_6_0_R0_en;
  wire [25:0] mem_6_0_W0_addr;
  wire  mem_6_0_W0_clk;
  wire [7:0] mem_6_0_W0_data;
  wire  mem_6_0_W0_en;
  wire  mem_6_0_W0_mask;
  wire [25:0] mem_6_1_R0_addr;
  wire  mem_6_1_R0_clk;
  wire [7:0] mem_6_1_R0_data;
  wire  mem_6_1_R0_en;
  wire [25:0] mem_6_1_W0_addr;
  wire  mem_6_1_W0_clk;
  wire [7:0] mem_6_1_W0_data;
  wire  mem_6_1_W0_en;
  wire  mem_6_1_W0_mask;
  wire [25:0] mem_6_2_R0_addr;
  wire  mem_6_2_R0_clk;
  wire [7:0] mem_6_2_R0_data;
  wire  mem_6_2_R0_en;
  wire [25:0] mem_6_2_W0_addr;
  wire  mem_6_2_W0_clk;
  wire [7:0] mem_6_2_W0_data;
  wire  mem_6_2_W0_en;
  wire  mem_6_2_W0_mask;
  wire [25:0] mem_6_3_R0_addr;
  wire  mem_6_3_R0_clk;
  wire [7:0] mem_6_3_R0_data;
  wire  mem_6_3_R0_en;
  wire [25:0] mem_6_3_W0_addr;
  wire  mem_6_3_W0_clk;
  wire [7:0] mem_6_3_W0_data;
  wire  mem_6_3_W0_en;
  wire  mem_6_3_W0_mask;
  wire [25:0] mem_6_4_R0_addr;
  wire  mem_6_4_R0_clk;
  wire [7:0] mem_6_4_R0_data;
  wire  mem_6_4_R0_en;
  wire [25:0] mem_6_4_W0_addr;
  wire  mem_6_4_W0_clk;
  wire [7:0] mem_6_4_W0_data;
  wire  mem_6_4_W0_en;
  wire  mem_6_4_W0_mask;
  wire [25:0] mem_6_5_R0_addr;
  wire  mem_6_5_R0_clk;
  wire [7:0] mem_6_5_R0_data;
  wire  mem_6_5_R0_en;
  wire [25:0] mem_6_5_W0_addr;
  wire  mem_6_5_W0_clk;
  wire [7:0] mem_6_5_W0_data;
  wire  mem_6_5_W0_en;
  wire  mem_6_5_W0_mask;
  wire [25:0] mem_6_6_R0_addr;
  wire  mem_6_6_R0_clk;
  wire [7:0] mem_6_6_R0_data;
  wire  mem_6_6_R0_en;
  wire [25:0] mem_6_6_W0_addr;
  wire  mem_6_6_W0_clk;
  wire [7:0] mem_6_6_W0_data;
  wire  mem_6_6_W0_en;
  wire  mem_6_6_W0_mask;
  wire [25:0] mem_6_7_R0_addr;
  wire  mem_6_7_R0_clk;
  wire [7:0] mem_6_7_R0_data;
  wire  mem_6_7_R0_en;
  wire [25:0] mem_6_7_W0_addr;
  wire  mem_6_7_W0_clk;
  wire [7:0] mem_6_7_W0_data;
  wire  mem_6_7_W0_en;
  wire  mem_6_7_W0_mask;
  wire [25:0] mem_7_0_R0_addr;
  wire  mem_7_0_R0_clk;
  wire [7:0] mem_7_0_R0_data;
  wire  mem_7_0_R0_en;
  wire [25:0] mem_7_0_W0_addr;
  wire  mem_7_0_W0_clk;
  wire [7:0] mem_7_0_W0_data;
  wire  mem_7_0_W0_en;
  wire  mem_7_0_W0_mask;
  wire [25:0] mem_7_1_R0_addr;
  wire  mem_7_1_R0_clk;
  wire [7:0] mem_7_1_R0_data;
  wire  mem_7_1_R0_en;
  wire [25:0] mem_7_1_W0_addr;
  wire  mem_7_1_W0_clk;
  wire [7:0] mem_7_1_W0_data;
  wire  mem_7_1_W0_en;
  wire  mem_7_1_W0_mask;
  wire [25:0] mem_7_2_R0_addr;
  wire  mem_7_2_R0_clk;
  wire [7:0] mem_7_2_R0_data;
  wire  mem_7_2_R0_en;
  wire [25:0] mem_7_2_W0_addr;
  wire  mem_7_2_W0_clk;
  wire [7:0] mem_7_2_W0_data;
  wire  mem_7_2_W0_en;
  wire  mem_7_2_W0_mask;
  wire [25:0] mem_7_3_R0_addr;
  wire  mem_7_3_R0_clk;
  wire [7:0] mem_7_3_R0_data;
  wire  mem_7_3_R0_en;
  wire [25:0] mem_7_3_W0_addr;
  wire  mem_7_3_W0_clk;
  wire [7:0] mem_7_3_W0_data;
  wire  mem_7_3_W0_en;
  wire  mem_7_3_W0_mask;
  wire [25:0] mem_7_4_R0_addr;
  wire  mem_7_4_R0_clk;
  wire [7:0] mem_7_4_R0_data;
  wire  mem_7_4_R0_en;
  wire [25:0] mem_7_4_W0_addr;
  wire  mem_7_4_W0_clk;
  wire [7:0] mem_7_4_W0_data;
  wire  mem_7_4_W0_en;
  wire  mem_7_4_W0_mask;
  wire [25:0] mem_7_5_R0_addr;
  wire  mem_7_5_R0_clk;
  wire [7:0] mem_7_5_R0_data;
  wire  mem_7_5_R0_en;
  wire [25:0] mem_7_5_W0_addr;
  wire  mem_7_5_W0_clk;
  wire [7:0] mem_7_5_W0_data;
  wire  mem_7_5_W0_en;
  wire  mem_7_5_W0_mask;
  wire [25:0] mem_7_6_R0_addr;
  wire  mem_7_6_R0_clk;
  wire [7:0] mem_7_6_R0_data;
  wire  mem_7_6_R0_en;
  wire [25:0] mem_7_6_W0_addr;
  wire  mem_7_6_W0_clk;
  wire [7:0] mem_7_6_W0_data;
  wire  mem_7_6_W0_en;
  wire  mem_7_6_W0_mask;
  wire [25:0] mem_7_7_R0_addr;
  wire  mem_7_7_R0_clk;
  wire [7:0] mem_7_7_R0_data;
  wire  mem_7_7_R0_en;
  wire [25:0] mem_7_7_W0_addr;
  wire  mem_7_7_W0_clk;
  wire [7:0] mem_7_7_W0_data;
  wire  mem_7_7_W0_en;
  wire  mem_7_7_W0_mask;
  wire [25:0] mem_8_0_R0_addr;
  wire  mem_8_0_R0_clk;
  wire [7:0] mem_8_0_R0_data;
  wire  mem_8_0_R0_en;
  wire [25:0] mem_8_0_W0_addr;
  wire  mem_8_0_W0_clk;
  wire [7:0] mem_8_0_W0_data;
  wire  mem_8_0_W0_en;
  wire  mem_8_0_W0_mask;
  wire [25:0] mem_8_1_R0_addr;
  wire  mem_8_1_R0_clk;
  wire [7:0] mem_8_1_R0_data;
  wire  mem_8_1_R0_en;
  wire [25:0] mem_8_1_W0_addr;
  wire  mem_8_1_W0_clk;
  wire [7:0] mem_8_1_W0_data;
  wire  mem_8_1_W0_en;
  wire  mem_8_1_W0_mask;
  wire [25:0] mem_8_2_R0_addr;
  wire  mem_8_2_R0_clk;
  wire [7:0] mem_8_2_R0_data;
  wire  mem_8_2_R0_en;
  wire [25:0] mem_8_2_W0_addr;
  wire  mem_8_2_W0_clk;
  wire [7:0] mem_8_2_W0_data;
  wire  mem_8_2_W0_en;
  wire  mem_8_2_W0_mask;
  wire [25:0] mem_8_3_R0_addr;
  wire  mem_8_3_R0_clk;
  wire [7:0] mem_8_3_R0_data;
  wire  mem_8_3_R0_en;
  wire [25:0] mem_8_3_W0_addr;
  wire  mem_8_3_W0_clk;
  wire [7:0] mem_8_3_W0_data;
  wire  mem_8_3_W0_en;
  wire  mem_8_3_W0_mask;
  wire [25:0] mem_8_4_R0_addr;
  wire  mem_8_4_R0_clk;
  wire [7:0] mem_8_4_R0_data;
  wire  mem_8_4_R0_en;
  wire [25:0] mem_8_4_W0_addr;
  wire  mem_8_4_W0_clk;
  wire [7:0] mem_8_4_W0_data;
  wire  mem_8_4_W0_en;
  wire  mem_8_4_W0_mask;
  wire [25:0] mem_8_5_R0_addr;
  wire  mem_8_5_R0_clk;
  wire [7:0] mem_8_5_R0_data;
  wire  mem_8_5_R0_en;
  wire [25:0] mem_8_5_W0_addr;
  wire  mem_8_5_W0_clk;
  wire [7:0] mem_8_5_W0_data;
  wire  mem_8_5_W0_en;
  wire  mem_8_5_W0_mask;
  wire [25:0] mem_8_6_R0_addr;
  wire  mem_8_6_R0_clk;
  wire [7:0] mem_8_6_R0_data;
  wire  mem_8_6_R0_en;
  wire [25:0] mem_8_6_W0_addr;
  wire  mem_8_6_W0_clk;
  wire [7:0] mem_8_6_W0_data;
  wire  mem_8_6_W0_en;
  wire  mem_8_6_W0_mask;
  wire [25:0] mem_8_7_R0_addr;
  wire  mem_8_7_R0_clk;
  wire [7:0] mem_8_7_R0_data;
  wire  mem_8_7_R0_en;
  wire [25:0] mem_8_7_W0_addr;
  wire  mem_8_7_W0_clk;
  wire [7:0] mem_8_7_W0_data;
  wire  mem_8_7_W0_en;
  wire  mem_8_7_W0_mask;
  wire [25:0] mem_9_0_R0_addr;
  wire  mem_9_0_R0_clk;
  wire [7:0] mem_9_0_R0_data;
  wire  mem_9_0_R0_en;
  wire [25:0] mem_9_0_W0_addr;
  wire  mem_9_0_W0_clk;
  wire [7:0] mem_9_0_W0_data;
  wire  mem_9_0_W0_en;
  wire  mem_9_0_W0_mask;
  wire [25:0] mem_9_1_R0_addr;
  wire  mem_9_1_R0_clk;
  wire [7:0] mem_9_1_R0_data;
  wire  mem_9_1_R0_en;
  wire [25:0] mem_9_1_W0_addr;
  wire  mem_9_1_W0_clk;
  wire [7:0] mem_9_1_W0_data;
  wire  mem_9_1_W0_en;
  wire  mem_9_1_W0_mask;
  wire [25:0] mem_9_2_R0_addr;
  wire  mem_9_2_R0_clk;
  wire [7:0] mem_9_2_R0_data;
  wire  mem_9_2_R0_en;
  wire [25:0] mem_9_2_W0_addr;
  wire  mem_9_2_W0_clk;
  wire [7:0] mem_9_2_W0_data;
  wire  mem_9_2_W0_en;
  wire  mem_9_2_W0_mask;
  wire [25:0] mem_9_3_R0_addr;
  wire  mem_9_3_R0_clk;
  wire [7:0] mem_9_3_R0_data;
  wire  mem_9_3_R0_en;
  wire [25:0] mem_9_3_W0_addr;
  wire  mem_9_3_W0_clk;
  wire [7:0] mem_9_3_W0_data;
  wire  mem_9_3_W0_en;
  wire  mem_9_3_W0_mask;
  wire [25:0] mem_9_4_R0_addr;
  wire  mem_9_4_R0_clk;
  wire [7:0] mem_9_4_R0_data;
  wire  mem_9_4_R0_en;
  wire [25:0] mem_9_4_W0_addr;
  wire  mem_9_4_W0_clk;
  wire [7:0] mem_9_4_W0_data;
  wire  mem_9_4_W0_en;
  wire  mem_9_4_W0_mask;
  wire [25:0] mem_9_5_R0_addr;
  wire  mem_9_5_R0_clk;
  wire [7:0] mem_9_5_R0_data;
  wire  mem_9_5_R0_en;
  wire [25:0] mem_9_5_W0_addr;
  wire  mem_9_5_W0_clk;
  wire [7:0] mem_9_5_W0_data;
  wire  mem_9_5_W0_en;
  wire  mem_9_5_W0_mask;
  wire [25:0] mem_9_6_R0_addr;
  wire  mem_9_6_R0_clk;
  wire [7:0] mem_9_6_R0_data;
  wire  mem_9_6_R0_en;
  wire [25:0] mem_9_6_W0_addr;
  wire  mem_9_6_W0_clk;
  wire [7:0] mem_9_6_W0_data;
  wire  mem_9_6_W0_en;
  wire  mem_9_6_W0_mask;
  wire [25:0] mem_9_7_R0_addr;
  wire  mem_9_7_R0_clk;
  wire [7:0] mem_9_7_R0_data;
  wire  mem_9_7_R0_en;
  wire [25:0] mem_9_7_W0_addr;
  wire  mem_9_7_W0_clk;
  wire [7:0] mem_9_7_W0_data;
  wire  mem_9_7_W0_en;
  wire  mem_9_7_W0_mask;
  wire [25:0] mem_10_0_R0_addr;
  wire  mem_10_0_R0_clk;
  wire [7:0] mem_10_0_R0_data;
  wire  mem_10_0_R0_en;
  wire [25:0] mem_10_0_W0_addr;
  wire  mem_10_0_W0_clk;
  wire [7:0] mem_10_0_W0_data;
  wire  mem_10_0_W0_en;
  wire  mem_10_0_W0_mask;
  wire [25:0] mem_10_1_R0_addr;
  wire  mem_10_1_R0_clk;
  wire [7:0] mem_10_1_R0_data;
  wire  mem_10_1_R0_en;
  wire [25:0] mem_10_1_W0_addr;
  wire  mem_10_1_W0_clk;
  wire [7:0] mem_10_1_W0_data;
  wire  mem_10_1_W0_en;
  wire  mem_10_1_W0_mask;
  wire [25:0] mem_10_2_R0_addr;
  wire  mem_10_2_R0_clk;
  wire [7:0] mem_10_2_R0_data;
  wire  mem_10_2_R0_en;
  wire [25:0] mem_10_2_W0_addr;
  wire  mem_10_2_W0_clk;
  wire [7:0] mem_10_2_W0_data;
  wire  mem_10_2_W0_en;
  wire  mem_10_2_W0_mask;
  wire [25:0] mem_10_3_R0_addr;
  wire  mem_10_3_R0_clk;
  wire [7:0] mem_10_3_R0_data;
  wire  mem_10_3_R0_en;
  wire [25:0] mem_10_3_W0_addr;
  wire  mem_10_3_W0_clk;
  wire [7:0] mem_10_3_W0_data;
  wire  mem_10_3_W0_en;
  wire  mem_10_3_W0_mask;
  wire [25:0] mem_10_4_R0_addr;
  wire  mem_10_4_R0_clk;
  wire [7:0] mem_10_4_R0_data;
  wire  mem_10_4_R0_en;
  wire [25:0] mem_10_4_W0_addr;
  wire  mem_10_4_W0_clk;
  wire [7:0] mem_10_4_W0_data;
  wire  mem_10_4_W0_en;
  wire  mem_10_4_W0_mask;
  wire [25:0] mem_10_5_R0_addr;
  wire  mem_10_5_R0_clk;
  wire [7:0] mem_10_5_R0_data;
  wire  mem_10_5_R0_en;
  wire [25:0] mem_10_5_W0_addr;
  wire  mem_10_5_W0_clk;
  wire [7:0] mem_10_5_W0_data;
  wire  mem_10_5_W0_en;
  wire  mem_10_5_W0_mask;
  wire [25:0] mem_10_6_R0_addr;
  wire  mem_10_6_R0_clk;
  wire [7:0] mem_10_6_R0_data;
  wire  mem_10_6_R0_en;
  wire [25:0] mem_10_6_W0_addr;
  wire  mem_10_6_W0_clk;
  wire [7:0] mem_10_6_W0_data;
  wire  mem_10_6_W0_en;
  wire  mem_10_6_W0_mask;
  wire [25:0] mem_10_7_R0_addr;
  wire  mem_10_7_R0_clk;
  wire [7:0] mem_10_7_R0_data;
  wire  mem_10_7_R0_en;
  wire [25:0] mem_10_7_W0_addr;
  wire  mem_10_7_W0_clk;
  wire [7:0] mem_10_7_W0_data;
  wire  mem_10_7_W0_en;
  wire  mem_10_7_W0_mask;
  wire [25:0] mem_11_0_R0_addr;
  wire  mem_11_0_R0_clk;
  wire [7:0] mem_11_0_R0_data;
  wire  mem_11_0_R0_en;
  wire [25:0] mem_11_0_W0_addr;
  wire  mem_11_0_W0_clk;
  wire [7:0] mem_11_0_W0_data;
  wire  mem_11_0_W0_en;
  wire  mem_11_0_W0_mask;
  wire [25:0] mem_11_1_R0_addr;
  wire  mem_11_1_R0_clk;
  wire [7:0] mem_11_1_R0_data;
  wire  mem_11_1_R0_en;
  wire [25:0] mem_11_1_W0_addr;
  wire  mem_11_1_W0_clk;
  wire [7:0] mem_11_1_W0_data;
  wire  mem_11_1_W0_en;
  wire  mem_11_1_W0_mask;
  wire [25:0] mem_11_2_R0_addr;
  wire  mem_11_2_R0_clk;
  wire [7:0] mem_11_2_R0_data;
  wire  mem_11_2_R0_en;
  wire [25:0] mem_11_2_W0_addr;
  wire  mem_11_2_W0_clk;
  wire [7:0] mem_11_2_W0_data;
  wire  mem_11_2_W0_en;
  wire  mem_11_2_W0_mask;
  wire [25:0] mem_11_3_R0_addr;
  wire  mem_11_3_R0_clk;
  wire [7:0] mem_11_3_R0_data;
  wire  mem_11_3_R0_en;
  wire [25:0] mem_11_3_W0_addr;
  wire  mem_11_3_W0_clk;
  wire [7:0] mem_11_3_W0_data;
  wire  mem_11_3_W0_en;
  wire  mem_11_3_W0_mask;
  wire [25:0] mem_11_4_R0_addr;
  wire  mem_11_4_R0_clk;
  wire [7:0] mem_11_4_R0_data;
  wire  mem_11_4_R0_en;
  wire [25:0] mem_11_4_W0_addr;
  wire  mem_11_4_W0_clk;
  wire [7:0] mem_11_4_W0_data;
  wire  mem_11_4_W0_en;
  wire  mem_11_4_W0_mask;
  wire [25:0] mem_11_5_R0_addr;
  wire  mem_11_5_R0_clk;
  wire [7:0] mem_11_5_R0_data;
  wire  mem_11_5_R0_en;
  wire [25:0] mem_11_5_W0_addr;
  wire  mem_11_5_W0_clk;
  wire [7:0] mem_11_5_W0_data;
  wire  mem_11_5_W0_en;
  wire  mem_11_5_W0_mask;
  wire [25:0] mem_11_6_R0_addr;
  wire  mem_11_6_R0_clk;
  wire [7:0] mem_11_6_R0_data;
  wire  mem_11_6_R0_en;
  wire [25:0] mem_11_6_W0_addr;
  wire  mem_11_6_W0_clk;
  wire [7:0] mem_11_6_W0_data;
  wire  mem_11_6_W0_en;
  wire  mem_11_6_W0_mask;
  wire [25:0] mem_11_7_R0_addr;
  wire  mem_11_7_R0_clk;
  wire [7:0] mem_11_7_R0_data;
  wire  mem_11_7_R0_en;
  wire [25:0] mem_11_7_W0_addr;
  wire  mem_11_7_W0_clk;
  wire [7:0] mem_11_7_W0_data;
  wire  mem_11_7_W0_en;
  wire  mem_11_7_W0_mask;
  wire [25:0] mem_12_0_R0_addr;
  wire  mem_12_0_R0_clk;
  wire [7:0] mem_12_0_R0_data;
  wire  mem_12_0_R0_en;
  wire [25:0] mem_12_0_W0_addr;
  wire  mem_12_0_W0_clk;
  wire [7:0] mem_12_0_W0_data;
  wire  mem_12_0_W0_en;
  wire  mem_12_0_W0_mask;
  wire [25:0] mem_12_1_R0_addr;
  wire  mem_12_1_R0_clk;
  wire [7:0] mem_12_1_R0_data;
  wire  mem_12_1_R0_en;
  wire [25:0] mem_12_1_W0_addr;
  wire  mem_12_1_W0_clk;
  wire [7:0] mem_12_1_W0_data;
  wire  mem_12_1_W0_en;
  wire  mem_12_1_W0_mask;
  wire [25:0] mem_12_2_R0_addr;
  wire  mem_12_2_R0_clk;
  wire [7:0] mem_12_2_R0_data;
  wire  mem_12_2_R0_en;
  wire [25:0] mem_12_2_W0_addr;
  wire  mem_12_2_W0_clk;
  wire [7:0] mem_12_2_W0_data;
  wire  mem_12_2_W0_en;
  wire  mem_12_2_W0_mask;
  wire [25:0] mem_12_3_R0_addr;
  wire  mem_12_3_R0_clk;
  wire [7:0] mem_12_3_R0_data;
  wire  mem_12_3_R0_en;
  wire [25:0] mem_12_3_W0_addr;
  wire  mem_12_3_W0_clk;
  wire [7:0] mem_12_3_W0_data;
  wire  mem_12_3_W0_en;
  wire  mem_12_3_W0_mask;
  wire [25:0] mem_12_4_R0_addr;
  wire  mem_12_4_R0_clk;
  wire [7:0] mem_12_4_R0_data;
  wire  mem_12_4_R0_en;
  wire [25:0] mem_12_4_W0_addr;
  wire  mem_12_4_W0_clk;
  wire [7:0] mem_12_4_W0_data;
  wire  mem_12_4_W0_en;
  wire  mem_12_4_W0_mask;
  wire [25:0] mem_12_5_R0_addr;
  wire  mem_12_5_R0_clk;
  wire [7:0] mem_12_5_R0_data;
  wire  mem_12_5_R0_en;
  wire [25:0] mem_12_5_W0_addr;
  wire  mem_12_5_W0_clk;
  wire [7:0] mem_12_5_W0_data;
  wire  mem_12_5_W0_en;
  wire  mem_12_5_W0_mask;
  wire [25:0] mem_12_6_R0_addr;
  wire  mem_12_6_R0_clk;
  wire [7:0] mem_12_6_R0_data;
  wire  mem_12_6_R0_en;
  wire [25:0] mem_12_6_W0_addr;
  wire  mem_12_6_W0_clk;
  wire [7:0] mem_12_6_W0_data;
  wire  mem_12_6_W0_en;
  wire  mem_12_6_W0_mask;
  wire [25:0] mem_12_7_R0_addr;
  wire  mem_12_7_R0_clk;
  wire [7:0] mem_12_7_R0_data;
  wire  mem_12_7_R0_en;
  wire [25:0] mem_12_7_W0_addr;
  wire  mem_12_7_W0_clk;
  wire [7:0] mem_12_7_W0_data;
  wire  mem_12_7_W0_en;
  wire  mem_12_7_W0_mask;
  wire [25:0] mem_13_0_R0_addr;
  wire  mem_13_0_R0_clk;
  wire [7:0] mem_13_0_R0_data;
  wire  mem_13_0_R0_en;
  wire [25:0] mem_13_0_W0_addr;
  wire  mem_13_0_W0_clk;
  wire [7:0] mem_13_0_W0_data;
  wire  mem_13_0_W0_en;
  wire  mem_13_0_W0_mask;
  wire [25:0] mem_13_1_R0_addr;
  wire  mem_13_1_R0_clk;
  wire [7:0] mem_13_1_R0_data;
  wire  mem_13_1_R0_en;
  wire [25:0] mem_13_1_W0_addr;
  wire  mem_13_1_W0_clk;
  wire [7:0] mem_13_1_W0_data;
  wire  mem_13_1_W0_en;
  wire  mem_13_1_W0_mask;
  wire [25:0] mem_13_2_R0_addr;
  wire  mem_13_2_R0_clk;
  wire [7:0] mem_13_2_R0_data;
  wire  mem_13_2_R0_en;
  wire [25:0] mem_13_2_W0_addr;
  wire  mem_13_2_W0_clk;
  wire [7:0] mem_13_2_W0_data;
  wire  mem_13_2_W0_en;
  wire  mem_13_2_W0_mask;
  wire [25:0] mem_13_3_R0_addr;
  wire  mem_13_3_R0_clk;
  wire [7:0] mem_13_3_R0_data;
  wire  mem_13_3_R0_en;
  wire [25:0] mem_13_3_W0_addr;
  wire  mem_13_3_W0_clk;
  wire [7:0] mem_13_3_W0_data;
  wire  mem_13_3_W0_en;
  wire  mem_13_3_W0_mask;
  wire [25:0] mem_13_4_R0_addr;
  wire  mem_13_4_R0_clk;
  wire [7:0] mem_13_4_R0_data;
  wire  mem_13_4_R0_en;
  wire [25:0] mem_13_4_W0_addr;
  wire  mem_13_4_W0_clk;
  wire [7:0] mem_13_4_W0_data;
  wire  mem_13_4_W0_en;
  wire  mem_13_4_W0_mask;
  wire [25:0] mem_13_5_R0_addr;
  wire  mem_13_5_R0_clk;
  wire [7:0] mem_13_5_R0_data;
  wire  mem_13_5_R0_en;
  wire [25:0] mem_13_5_W0_addr;
  wire  mem_13_5_W0_clk;
  wire [7:0] mem_13_5_W0_data;
  wire  mem_13_5_W0_en;
  wire  mem_13_5_W0_mask;
  wire [25:0] mem_13_6_R0_addr;
  wire  mem_13_6_R0_clk;
  wire [7:0] mem_13_6_R0_data;
  wire  mem_13_6_R0_en;
  wire [25:0] mem_13_6_W0_addr;
  wire  mem_13_6_W0_clk;
  wire [7:0] mem_13_6_W0_data;
  wire  mem_13_6_W0_en;
  wire  mem_13_6_W0_mask;
  wire [25:0] mem_13_7_R0_addr;
  wire  mem_13_7_R0_clk;
  wire [7:0] mem_13_7_R0_data;
  wire  mem_13_7_R0_en;
  wire [25:0] mem_13_7_W0_addr;
  wire  mem_13_7_W0_clk;
  wire [7:0] mem_13_7_W0_data;
  wire  mem_13_7_W0_en;
  wire  mem_13_7_W0_mask;
  wire [25:0] mem_14_0_R0_addr;
  wire  mem_14_0_R0_clk;
  wire [7:0] mem_14_0_R0_data;
  wire  mem_14_0_R0_en;
  wire [25:0] mem_14_0_W0_addr;
  wire  mem_14_0_W0_clk;
  wire [7:0] mem_14_0_W0_data;
  wire  mem_14_0_W0_en;
  wire  mem_14_0_W0_mask;
  wire [25:0] mem_14_1_R0_addr;
  wire  mem_14_1_R0_clk;
  wire [7:0] mem_14_1_R0_data;
  wire  mem_14_1_R0_en;
  wire [25:0] mem_14_1_W0_addr;
  wire  mem_14_1_W0_clk;
  wire [7:0] mem_14_1_W0_data;
  wire  mem_14_1_W0_en;
  wire  mem_14_1_W0_mask;
  wire [25:0] mem_14_2_R0_addr;
  wire  mem_14_2_R0_clk;
  wire [7:0] mem_14_2_R0_data;
  wire  mem_14_2_R0_en;
  wire [25:0] mem_14_2_W0_addr;
  wire  mem_14_2_W0_clk;
  wire [7:0] mem_14_2_W0_data;
  wire  mem_14_2_W0_en;
  wire  mem_14_2_W0_mask;
  wire [25:0] mem_14_3_R0_addr;
  wire  mem_14_3_R0_clk;
  wire [7:0] mem_14_3_R0_data;
  wire  mem_14_3_R0_en;
  wire [25:0] mem_14_3_W0_addr;
  wire  mem_14_3_W0_clk;
  wire [7:0] mem_14_3_W0_data;
  wire  mem_14_3_W0_en;
  wire  mem_14_3_W0_mask;
  wire [25:0] mem_14_4_R0_addr;
  wire  mem_14_4_R0_clk;
  wire [7:0] mem_14_4_R0_data;
  wire  mem_14_4_R0_en;
  wire [25:0] mem_14_4_W0_addr;
  wire  mem_14_4_W0_clk;
  wire [7:0] mem_14_4_W0_data;
  wire  mem_14_4_W0_en;
  wire  mem_14_4_W0_mask;
  wire [25:0] mem_14_5_R0_addr;
  wire  mem_14_5_R0_clk;
  wire [7:0] mem_14_5_R0_data;
  wire  mem_14_5_R0_en;
  wire [25:0] mem_14_5_W0_addr;
  wire  mem_14_5_W0_clk;
  wire [7:0] mem_14_5_W0_data;
  wire  mem_14_5_W0_en;
  wire  mem_14_5_W0_mask;
  wire [25:0] mem_14_6_R0_addr;
  wire  mem_14_6_R0_clk;
  wire [7:0] mem_14_6_R0_data;
  wire  mem_14_6_R0_en;
  wire [25:0] mem_14_6_W0_addr;
  wire  mem_14_6_W0_clk;
  wire [7:0] mem_14_6_W0_data;
  wire  mem_14_6_W0_en;
  wire  mem_14_6_W0_mask;
  wire [25:0] mem_14_7_R0_addr;
  wire  mem_14_7_R0_clk;
  wire [7:0] mem_14_7_R0_data;
  wire  mem_14_7_R0_en;
  wire [25:0] mem_14_7_W0_addr;
  wire  mem_14_7_W0_clk;
  wire [7:0] mem_14_7_W0_data;
  wire  mem_14_7_W0_en;
  wire  mem_14_7_W0_mask;
  wire [25:0] mem_15_0_R0_addr;
  wire  mem_15_0_R0_clk;
  wire [7:0] mem_15_0_R0_data;
  wire  mem_15_0_R0_en;
  wire [25:0] mem_15_0_W0_addr;
  wire  mem_15_0_W0_clk;
  wire [7:0] mem_15_0_W0_data;
  wire  mem_15_0_W0_en;
  wire  mem_15_0_W0_mask;
  wire [25:0] mem_15_1_R0_addr;
  wire  mem_15_1_R0_clk;
  wire [7:0] mem_15_1_R0_data;
  wire  mem_15_1_R0_en;
  wire [25:0] mem_15_1_W0_addr;
  wire  mem_15_1_W0_clk;
  wire [7:0] mem_15_1_W0_data;
  wire  mem_15_1_W0_en;
  wire  mem_15_1_W0_mask;
  wire [25:0] mem_15_2_R0_addr;
  wire  mem_15_2_R0_clk;
  wire [7:0] mem_15_2_R0_data;
  wire  mem_15_2_R0_en;
  wire [25:0] mem_15_2_W0_addr;
  wire  mem_15_2_W0_clk;
  wire [7:0] mem_15_2_W0_data;
  wire  mem_15_2_W0_en;
  wire  mem_15_2_W0_mask;
  wire [25:0] mem_15_3_R0_addr;
  wire  mem_15_3_R0_clk;
  wire [7:0] mem_15_3_R0_data;
  wire  mem_15_3_R0_en;
  wire [25:0] mem_15_3_W0_addr;
  wire  mem_15_3_W0_clk;
  wire [7:0] mem_15_3_W0_data;
  wire  mem_15_3_W0_en;
  wire  mem_15_3_W0_mask;
  wire [25:0] mem_15_4_R0_addr;
  wire  mem_15_4_R0_clk;
  wire [7:0] mem_15_4_R0_data;
  wire  mem_15_4_R0_en;
  wire [25:0] mem_15_4_W0_addr;
  wire  mem_15_4_W0_clk;
  wire [7:0] mem_15_4_W0_data;
  wire  mem_15_4_W0_en;
  wire  mem_15_4_W0_mask;
  wire [25:0] mem_15_5_R0_addr;
  wire  mem_15_5_R0_clk;
  wire [7:0] mem_15_5_R0_data;
  wire  mem_15_5_R0_en;
  wire [25:0] mem_15_5_W0_addr;
  wire  mem_15_5_W0_clk;
  wire [7:0] mem_15_5_W0_data;
  wire  mem_15_5_W0_en;
  wire  mem_15_5_W0_mask;
  wire [25:0] mem_15_6_R0_addr;
  wire  mem_15_6_R0_clk;
  wire [7:0] mem_15_6_R0_data;
  wire  mem_15_6_R0_en;
  wire [25:0] mem_15_6_W0_addr;
  wire  mem_15_6_W0_clk;
  wire [7:0] mem_15_6_W0_data;
  wire  mem_15_6_W0_en;
  wire  mem_15_6_W0_mask;
  wire [25:0] mem_15_7_R0_addr;
  wire  mem_15_7_R0_clk;
  wire [7:0] mem_15_7_R0_data;
  wire  mem_15_7_R0_en;
  wire [25:0] mem_15_7_W0_addr;
  wire  mem_15_7_W0_clk;
  wire [7:0] mem_15_7_W0_data;
  wire  mem_15_7_W0_en;
  wire  mem_15_7_W0_mask;
  wire [25:0] mem_16_0_R0_addr;
  wire  mem_16_0_R0_clk;
  wire [7:0] mem_16_0_R0_data;
  wire  mem_16_0_R0_en;
  wire [25:0] mem_16_0_W0_addr;
  wire  mem_16_0_W0_clk;
  wire [7:0] mem_16_0_W0_data;
  wire  mem_16_0_W0_en;
  wire  mem_16_0_W0_mask;
  wire [25:0] mem_16_1_R0_addr;
  wire  mem_16_1_R0_clk;
  wire [7:0] mem_16_1_R0_data;
  wire  mem_16_1_R0_en;
  wire [25:0] mem_16_1_W0_addr;
  wire  mem_16_1_W0_clk;
  wire [7:0] mem_16_1_W0_data;
  wire  mem_16_1_W0_en;
  wire  mem_16_1_W0_mask;
  wire [25:0] mem_16_2_R0_addr;
  wire  mem_16_2_R0_clk;
  wire [7:0] mem_16_2_R0_data;
  wire  mem_16_2_R0_en;
  wire [25:0] mem_16_2_W0_addr;
  wire  mem_16_2_W0_clk;
  wire [7:0] mem_16_2_W0_data;
  wire  mem_16_2_W0_en;
  wire  mem_16_2_W0_mask;
  wire [25:0] mem_16_3_R0_addr;
  wire  mem_16_3_R0_clk;
  wire [7:0] mem_16_3_R0_data;
  wire  mem_16_3_R0_en;
  wire [25:0] mem_16_3_W0_addr;
  wire  mem_16_3_W0_clk;
  wire [7:0] mem_16_3_W0_data;
  wire  mem_16_3_W0_en;
  wire  mem_16_3_W0_mask;
  wire [25:0] mem_16_4_R0_addr;
  wire  mem_16_4_R0_clk;
  wire [7:0] mem_16_4_R0_data;
  wire  mem_16_4_R0_en;
  wire [25:0] mem_16_4_W0_addr;
  wire  mem_16_4_W0_clk;
  wire [7:0] mem_16_4_W0_data;
  wire  mem_16_4_W0_en;
  wire  mem_16_4_W0_mask;
  wire [25:0] mem_16_5_R0_addr;
  wire  mem_16_5_R0_clk;
  wire [7:0] mem_16_5_R0_data;
  wire  mem_16_5_R0_en;
  wire [25:0] mem_16_5_W0_addr;
  wire  mem_16_5_W0_clk;
  wire [7:0] mem_16_5_W0_data;
  wire  mem_16_5_W0_en;
  wire  mem_16_5_W0_mask;
  wire [25:0] mem_16_6_R0_addr;
  wire  mem_16_6_R0_clk;
  wire [7:0] mem_16_6_R0_data;
  wire  mem_16_6_R0_en;
  wire [25:0] mem_16_6_W0_addr;
  wire  mem_16_6_W0_clk;
  wire [7:0] mem_16_6_W0_data;
  wire  mem_16_6_W0_en;
  wire  mem_16_6_W0_mask;
  wire [25:0] mem_16_7_R0_addr;
  wire  mem_16_7_R0_clk;
  wire [7:0] mem_16_7_R0_data;
  wire  mem_16_7_R0_en;
  wire [25:0] mem_16_7_W0_addr;
  wire  mem_16_7_W0_clk;
  wire [7:0] mem_16_7_W0_data;
  wire  mem_16_7_W0_en;
  wire  mem_16_7_W0_mask;
  wire [25:0] mem_17_0_R0_addr;
  wire  mem_17_0_R0_clk;
  wire [7:0] mem_17_0_R0_data;
  wire  mem_17_0_R0_en;
  wire [25:0] mem_17_0_W0_addr;
  wire  mem_17_0_W0_clk;
  wire [7:0] mem_17_0_W0_data;
  wire  mem_17_0_W0_en;
  wire  mem_17_0_W0_mask;
  wire [25:0] mem_17_1_R0_addr;
  wire  mem_17_1_R0_clk;
  wire [7:0] mem_17_1_R0_data;
  wire  mem_17_1_R0_en;
  wire [25:0] mem_17_1_W0_addr;
  wire  mem_17_1_W0_clk;
  wire [7:0] mem_17_1_W0_data;
  wire  mem_17_1_W0_en;
  wire  mem_17_1_W0_mask;
  wire [25:0] mem_17_2_R0_addr;
  wire  mem_17_2_R0_clk;
  wire [7:0] mem_17_2_R0_data;
  wire  mem_17_2_R0_en;
  wire [25:0] mem_17_2_W0_addr;
  wire  mem_17_2_W0_clk;
  wire [7:0] mem_17_2_W0_data;
  wire  mem_17_2_W0_en;
  wire  mem_17_2_W0_mask;
  wire [25:0] mem_17_3_R0_addr;
  wire  mem_17_3_R0_clk;
  wire [7:0] mem_17_3_R0_data;
  wire  mem_17_3_R0_en;
  wire [25:0] mem_17_3_W0_addr;
  wire  mem_17_3_W0_clk;
  wire [7:0] mem_17_3_W0_data;
  wire  mem_17_3_W0_en;
  wire  mem_17_3_W0_mask;
  wire [25:0] mem_17_4_R0_addr;
  wire  mem_17_4_R0_clk;
  wire [7:0] mem_17_4_R0_data;
  wire  mem_17_4_R0_en;
  wire [25:0] mem_17_4_W0_addr;
  wire  mem_17_4_W0_clk;
  wire [7:0] mem_17_4_W0_data;
  wire  mem_17_4_W0_en;
  wire  mem_17_4_W0_mask;
  wire [25:0] mem_17_5_R0_addr;
  wire  mem_17_5_R0_clk;
  wire [7:0] mem_17_5_R0_data;
  wire  mem_17_5_R0_en;
  wire [25:0] mem_17_5_W0_addr;
  wire  mem_17_5_W0_clk;
  wire [7:0] mem_17_5_W0_data;
  wire  mem_17_5_W0_en;
  wire  mem_17_5_W0_mask;
  wire [25:0] mem_17_6_R0_addr;
  wire  mem_17_6_R0_clk;
  wire [7:0] mem_17_6_R0_data;
  wire  mem_17_6_R0_en;
  wire [25:0] mem_17_6_W0_addr;
  wire  mem_17_6_W0_clk;
  wire [7:0] mem_17_6_W0_data;
  wire  mem_17_6_W0_en;
  wire  mem_17_6_W0_mask;
  wire [25:0] mem_17_7_R0_addr;
  wire  mem_17_7_R0_clk;
  wire [7:0] mem_17_7_R0_data;
  wire  mem_17_7_R0_en;
  wire [25:0] mem_17_7_W0_addr;
  wire  mem_17_7_W0_clk;
  wire [7:0] mem_17_7_W0_data;
  wire  mem_17_7_W0_en;
  wire  mem_17_7_W0_mask;
  wire [25:0] mem_18_0_R0_addr;
  wire  mem_18_0_R0_clk;
  wire [7:0] mem_18_0_R0_data;
  wire  mem_18_0_R0_en;
  wire [25:0] mem_18_0_W0_addr;
  wire  mem_18_0_W0_clk;
  wire [7:0] mem_18_0_W0_data;
  wire  mem_18_0_W0_en;
  wire  mem_18_0_W0_mask;
  wire [25:0] mem_18_1_R0_addr;
  wire  mem_18_1_R0_clk;
  wire [7:0] mem_18_1_R0_data;
  wire  mem_18_1_R0_en;
  wire [25:0] mem_18_1_W0_addr;
  wire  mem_18_1_W0_clk;
  wire [7:0] mem_18_1_W0_data;
  wire  mem_18_1_W0_en;
  wire  mem_18_1_W0_mask;
  wire [25:0] mem_18_2_R0_addr;
  wire  mem_18_2_R0_clk;
  wire [7:0] mem_18_2_R0_data;
  wire  mem_18_2_R0_en;
  wire [25:0] mem_18_2_W0_addr;
  wire  mem_18_2_W0_clk;
  wire [7:0] mem_18_2_W0_data;
  wire  mem_18_2_W0_en;
  wire  mem_18_2_W0_mask;
  wire [25:0] mem_18_3_R0_addr;
  wire  mem_18_3_R0_clk;
  wire [7:0] mem_18_3_R0_data;
  wire  mem_18_3_R0_en;
  wire [25:0] mem_18_3_W0_addr;
  wire  mem_18_3_W0_clk;
  wire [7:0] mem_18_3_W0_data;
  wire  mem_18_3_W0_en;
  wire  mem_18_3_W0_mask;
  wire [25:0] mem_18_4_R0_addr;
  wire  mem_18_4_R0_clk;
  wire [7:0] mem_18_4_R0_data;
  wire  mem_18_4_R0_en;
  wire [25:0] mem_18_4_W0_addr;
  wire  mem_18_4_W0_clk;
  wire [7:0] mem_18_4_W0_data;
  wire  mem_18_4_W0_en;
  wire  mem_18_4_W0_mask;
  wire [25:0] mem_18_5_R0_addr;
  wire  mem_18_5_R0_clk;
  wire [7:0] mem_18_5_R0_data;
  wire  mem_18_5_R0_en;
  wire [25:0] mem_18_5_W0_addr;
  wire  mem_18_5_W0_clk;
  wire [7:0] mem_18_5_W0_data;
  wire  mem_18_5_W0_en;
  wire  mem_18_5_W0_mask;
  wire [25:0] mem_18_6_R0_addr;
  wire  mem_18_6_R0_clk;
  wire [7:0] mem_18_6_R0_data;
  wire  mem_18_6_R0_en;
  wire [25:0] mem_18_6_W0_addr;
  wire  mem_18_6_W0_clk;
  wire [7:0] mem_18_6_W0_data;
  wire  mem_18_6_W0_en;
  wire  mem_18_6_W0_mask;
  wire [25:0] mem_18_7_R0_addr;
  wire  mem_18_7_R0_clk;
  wire [7:0] mem_18_7_R0_data;
  wire  mem_18_7_R0_en;
  wire [25:0] mem_18_7_W0_addr;
  wire  mem_18_7_W0_clk;
  wire [7:0] mem_18_7_W0_data;
  wire  mem_18_7_W0_en;
  wire  mem_18_7_W0_mask;
  wire [25:0] mem_19_0_R0_addr;
  wire  mem_19_0_R0_clk;
  wire [7:0] mem_19_0_R0_data;
  wire  mem_19_0_R0_en;
  wire [25:0] mem_19_0_W0_addr;
  wire  mem_19_0_W0_clk;
  wire [7:0] mem_19_0_W0_data;
  wire  mem_19_0_W0_en;
  wire  mem_19_0_W0_mask;
  wire [25:0] mem_19_1_R0_addr;
  wire  mem_19_1_R0_clk;
  wire [7:0] mem_19_1_R0_data;
  wire  mem_19_1_R0_en;
  wire [25:0] mem_19_1_W0_addr;
  wire  mem_19_1_W0_clk;
  wire [7:0] mem_19_1_W0_data;
  wire  mem_19_1_W0_en;
  wire  mem_19_1_W0_mask;
  wire [25:0] mem_19_2_R0_addr;
  wire  mem_19_2_R0_clk;
  wire [7:0] mem_19_2_R0_data;
  wire  mem_19_2_R0_en;
  wire [25:0] mem_19_2_W0_addr;
  wire  mem_19_2_W0_clk;
  wire [7:0] mem_19_2_W0_data;
  wire  mem_19_2_W0_en;
  wire  mem_19_2_W0_mask;
  wire [25:0] mem_19_3_R0_addr;
  wire  mem_19_3_R0_clk;
  wire [7:0] mem_19_3_R0_data;
  wire  mem_19_3_R0_en;
  wire [25:0] mem_19_3_W0_addr;
  wire  mem_19_3_W0_clk;
  wire [7:0] mem_19_3_W0_data;
  wire  mem_19_3_W0_en;
  wire  mem_19_3_W0_mask;
  wire [25:0] mem_19_4_R0_addr;
  wire  mem_19_4_R0_clk;
  wire [7:0] mem_19_4_R0_data;
  wire  mem_19_4_R0_en;
  wire [25:0] mem_19_4_W0_addr;
  wire  mem_19_4_W0_clk;
  wire [7:0] mem_19_4_W0_data;
  wire  mem_19_4_W0_en;
  wire  mem_19_4_W0_mask;
  wire [25:0] mem_19_5_R0_addr;
  wire  mem_19_5_R0_clk;
  wire [7:0] mem_19_5_R0_data;
  wire  mem_19_5_R0_en;
  wire [25:0] mem_19_5_W0_addr;
  wire  mem_19_5_W0_clk;
  wire [7:0] mem_19_5_W0_data;
  wire  mem_19_5_W0_en;
  wire  mem_19_5_W0_mask;
  wire [25:0] mem_19_6_R0_addr;
  wire  mem_19_6_R0_clk;
  wire [7:0] mem_19_6_R0_data;
  wire  mem_19_6_R0_en;
  wire [25:0] mem_19_6_W0_addr;
  wire  mem_19_6_W0_clk;
  wire [7:0] mem_19_6_W0_data;
  wire  mem_19_6_W0_en;
  wire  mem_19_6_W0_mask;
  wire [25:0] mem_19_7_R0_addr;
  wire  mem_19_7_R0_clk;
  wire [7:0] mem_19_7_R0_data;
  wire  mem_19_7_R0_en;
  wire [25:0] mem_19_7_W0_addr;
  wire  mem_19_7_W0_clk;
  wire [7:0] mem_19_7_W0_data;
  wire  mem_19_7_W0_en;
  wire  mem_19_7_W0_mask;
  wire [25:0] mem_20_0_R0_addr;
  wire  mem_20_0_R0_clk;
  wire [7:0] mem_20_0_R0_data;
  wire  mem_20_0_R0_en;
  wire [25:0] mem_20_0_W0_addr;
  wire  mem_20_0_W0_clk;
  wire [7:0] mem_20_0_W0_data;
  wire  mem_20_0_W0_en;
  wire  mem_20_0_W0_mask;
  wire [25:0] mem_20_1_R0_addr;
  wire  mem_20_1_R0_clk;
  wire [7:0] mem_20_1_R0_data;
  wire  mem_20_1_R0_en;
  wire [25:0] mem_20_1_W0_addr;
  wire  mem_20_1_W0_clk;
  wire [7:0] mem_20_1_W0_data;
  wire  mem_20_1_W0_en;
  wire  mem_20_1_W0_mask;
  wire [25:0] mem_20_2_R0_addr;
  wire  mem_20_2_R0_clk;
  wire [7:0] mem_20_2_R0_data;
  wire  mem_20_2_R0_en;
  wire [25:0] mem_20_2_W0_addr;
  wire  mem_20_2_W0_clk;
  wire [7:0] mem_20_2_W0_data;
  wire  mem_20_2_W0_en;
  wire  mem_20_2_W0_mask;
  wire [25:0] mem_20_3_R0_addr;
  wire  mem_20_3_R0_clk;
  wire [7:0] mem_20_3_R0_data;
  wire  mem_20_3_R0_en;
  wire [25:0] mem_20_3_W0_addr;
  wire  mem_20_3_W0_clk;
  wire [7:0] mem_20_3_W0_data;
  wire  mem_20_3_W0_en;
  wire  mem_20_3_W0_mask;
  wire [25:0] mem_20_4_R0_addr;
  wire  mem_20_4_R0_clk;
  wire [7:0] mem_20_4_R0_data;
  wire  mem_20_4_R0_en;
  wire [25:0] mem_20_4_W0_addr;
  wire  mem_20_4_W0_clk;
  wire [7:0] mem_20_4_W0_data;
  wire  mem_20_4_W0_en;
  wire  mem_20_4_W0_mask;
  wire [25:0] mem_20_5_R0_addr;
  wire  mem_20_5_R0_clk;
  wire [7:0] mem_20_5_R0_data;
  wire  mem_20_5_R0_en;
  wire [25:0] mem_20_5_W0_addr;
  wire  mem_20_5_W0_clk;
  wire [7:0] mem_20_5_W0_data;
  wire  mem_20_5_W0_en;
  wire  mem_20_5_W0_mask;
  wire [25:0] mem_20_6_R0_addr;
  wire  mem_20_6_R0_clk;
  wire [7:0] mem_20_6_R0_data;
  wire  mem_20_6_R0_en;
  wire [25:0] mem_20_6_W0_addr;
  wire  mem_20_6_W0_clk;
  wire [7:0] mem_20_6_W0_data;
  wire  mem_20_6_W0_en;
  wire  mem_20_6_W0_mask;
  wire [25:0] mem_20_7_R0_addr;
  wire  mem_20_7_R0_clk;
  wire [7:0] mem_20_7_R0_data;
  wire  mem_20_7_R0_en;
  wire [25:0] mem_20_7_W0_addr;
  wire  mem_20_7_W0_clk;
  wire [7:0] mem_20_7_W0_data;
  wire  mem_20_7_W0_en;
  wire  mem_20_7_W0_mask;
  wire [25:0] mem_21_0_R0_addr;
  wire  mem_21_0_R0_clk;
  wire [7:0] mem_21_0_R0_data;
  wire  mem_21_0_R0_en;
  wire [25:0] mem_21_0_W0_addr;
  wire  mem_21_0_W0_clk;
  wire [7:0] mem_21_0_W0_data;
  wire  mem_21_0_W0_en;
  wire  mem_21_0_W0_mask;
  wire [25:0] mem_21_1_R0_addr;
  wire  mem_21_1_R0_clk;
  wire [7:0] mem_21_1_R0_data;
  wire  mem_21_1_R0_en;
  wire [25:0] mem_21_1_W0_addr;
  wire  mem_21_1_W0_clk;
  wire [7:0] mem_21_1_W0_data;
  wire  mem_21_1_W0_en;
  wire  mem_21_1_W0_mask;
  wire [25:0] mem_21_2_R0_addr;
  wire  mem_21_2_R0_clk;
  wire [7:0] mem_21_2_R0_data;
  wire  mem_21_2_R0_en;
  wire [25:0] mem_21_2_W0_addr;
  wire  mem_21_2_W0_clk;
  wire [7:0] mem_21_2_W0_data;
  wire  mem_21_2_W0_en;
  wire  mem_21_2_W0_mask;
  wire [25:0] mem_21_3_R0_addr;
  wire  mem_21_3_R0_clk;
  wire [7:0] mem_21_3_R0_data;
  wire  mem_21_3_R0_en;
  wire [25:0] mem_21_3_W0_addr;
  wire  mem_21_3_W0_clk;
  wire [7:0] mem_21_3_W0_data;
  wire  mem_21_3_W0_en;
  wire  mem_21_3_W0_mask;
  wire [25:0] mem_21_4_R0_addr;
  wire  mem_21_4_R0_clk;
  wire [7:0] mem_21_4_R0_data;
  wire  mem_21_4_R0_en;
  wire [25:0] mem_21_4_W0_addr;
  wire  mem_21_4_W0_clk;
  wire [7:0] mem_21_4_W0_data;
  wire  mem_21_4_W0_en;
  wire  mem_21_4_W0_mask;
  wire [25:0] mem_21_5_R0_addr;
  wire  mem_21_5_R0_clk;
  wire [7:0] mem_21_5_R0_data;
  wire  mem_21_5_R0_en;
  wire [25:0] mem_21_5_W0_addr;
  wire  mem_21_5_W0_clk;
  wire [7:0] mem_21_5_W0_data;
  wire  mem_21_5_W0_en;
  wire  mem_21_5_W0_mask;
  wire [25:0] mem_21_6_R0_addr;
  wire  mem_21_6_R0_clk;
  wire [7:0] mem_21_6_R0_data;
  wire  mem_21_6_R0_en;
  wire [25:0] mem_21_6_W0_addr;
  wire  mem_21_6_W0_clk;
  wire [7:0] mem_21_6_W0_data;
  wire  mem_21_6_W0_en;
  wire  mem_21_6_W0_mask;
  wire [25:0] mem_21_7_R0_addr;
  wire  mem_21_7_R0_clk;
  wire [7:0] mem_21_7_R0_data;
  wire  mem_21_7_R0_en;
  wire [25:0] mem_21_7_W0_addr;
  wire  mem_21_7_W0_clk;
  wire [7:0] mem_21_7_W0_data;
  wire  mem_21_7_W0_en;
  wire  mem_21_7_W0_mask;
  wire [25:0] mem_22_0_R0_addr;
  wire  mem_22_0_R0_clk;
  wire [7:0] mem_22_0_R0_data;
  wire  mem_22_0_R0_en;
  wire [25:0] mem_22_0_W0_addr;
  wire  mem_22_0_W0_clk;
  wire [7:0] mem_22_0_W0_data;
  wire  mem_22_0_W0_en;
  wire  mem_22_0_W0_mask;
  wire [25:0] mem_22_1_R0_addr;
  wire  mem_22_1_R0_clk;
  wire [7:0] mem_22_1_R0_data;
  wire  mem_22_1_R0_en;
  wire [25:0] mem_22_1_W0_addr;
  wire  mem_22_1_W0_clk;
  wire [7:0] mem_22_1_W0_data;
  wire  mem_22_1_W0_en;
  wire  mem_22_1_W0_mask;
  wire [25:0] mem_22_2_R0_addr;
  wire  mem_22_2_R0_clk;
  wire [7:0] mem_22_2_R0_data;
  wire  mem_22_2_R0_en;
  wire [25:0] mem_22_2_W0_addr;
  wire  mem_22_2_W0_clk;
  wire [7:0] mem_22_2_W0_data;
  wire  mem_22_2_W0_en;
  wire  mem_22_2_W0_mask;
  wire [25:0] mem_22_3_R0_addr;
  wire  mem_22_3_R0_clk;
  wire [7:0] mem_22_3_R0_data;
  wire  mem_22_3_R0_en;
  wire [25:0] mem_22_3_W0_addr;
  wire  mem_22_3_W0_clk;
  wire [7:0] mem_22_3_W0_data;
  wire  mem_22_3_W0_en;
  wire  mem_22_3_W0_mask;
  wire [25:0] mem_22_4_R0_addr;
  wire  mem_22_4_R0_clk;
  wire [7:0] mem_22_4_R0_data;
  wire  mem_22_4_R0_en;
  wire [25:0] mem_22_4_W0_addr;
  wire  mem_22_4_W0_clk;
  wire [7:0] mem_22_4_W0_data;
  wire  mem_22_4_W0_en;
  wire  mem_22_4_W0_mask;
  wire [25:0] mem_22_5_R0_addr;
  wire  mem_22_5_R0_clk;
  wire [7:0] mem_22_5_R0_data;
  wire  mem_22_5_R0_en;
  wire [25:0] mem_22_5_W0_addr;
  wire  mem_22_5_W0_clk;
  wire [7:0] mem_22_5_W0_data;
  wire  mem_22_5_W0_en;
  wire  mem_22_5_W0_mask;
  wire [25:0] mem_22_6_R0_addr;
  wire  mem_22_6_R0_clk;
  wire [7:0] mem_22_6_R0_data;
  wire  mem_22_6_R0_en;
  wire [25:0] mem_22_6_W0_addr;
  wire  mem_22_6_W0_clk;
  wire [7:0] mem_22_6_W0_data;
  wire  mem_22_6_W0_en;
  wire  mem_22_6_W0_mask;
  wire [25:0] mem_22_7_R0_addr;
  wire  mem_22_7_R0_clk;
  wire [7:0] mem_22_7_R0_data;
  wire  mem_22_7_R0_en;
  wire [25:0] mem_22_7_W0_addr;
  wire  mem_22_7_W0_clk;
  wire [7:0] mem_22_7_W0_data;
  wire  mem_22_7_W0_en;
  wire  mem_22_7_W0_mask;
  wire [25:0] mem_23_0_R0_addr;
  wire  mem_23_0_R0_clk;
  wire [7:0] mem_23_0_R0_data;
  wire  mem_23_0_R0_en;
  wire [25:0] mem_23_0_W0_addr;
  wire  mem_23_0_W0_clk;
  wire [7:0] mem_23_0_W0_data;
  wire  mem_23_0_W0_en;
  wire  mem_23_0_W0_mask;
  wire [25:0] mem_23_1_R0_addr;
  wire  mem_23_1_R0_clk;
  wire [7:0] mem_23_1_R0_data;
  wire  mem_23_1_R0_en;
  wire [25:0] mem_23_1_W0_addr;
  wire  mem_23_1_W0_clk;
  wire [7:0] mem_23_1_W0_data;
  wire  mem_23_1_W0_en;
  wire  mem_23_1_W0_mask;
  wire [25:0] mem_23_2_R0_addr;
  wire  mem_23_2_R0_clk;
  wire [7:0] mem_23_2_R0_data;
  wire  mem_23_2_R0_en;
  wire [25:0] mem_23_2_W0_addr;
  wire  mem_23_2_W0_clk;
  wire [7:0] mem_23_2_W0_data;
  wire  mem_23_2_W0_en;
  wire  mem_23_2_W0_mask;
  wire [25:0] mem_23_3_R0_addr;
  wire  mem_23_3_R0_clk;
  wire [7:0] mem_23_3_R0_data;
  wire  mem_23_3_R0_en;
  wire [25:0] mem_23_3_W0_addr;
  wire  mem_23_3_W0_clk;
  wire [7:0] mem_23_3_W0_data;
  wire  mem_23_3_W0_en;
  wire  mem_23_3_W0_mask;
  wire [25:0] mem_23_4_R0_addr;
  wire  mem_23_4_R0_clk;
  wire [7:0] mem_23_4_R0_data;
  wire  mem_23_4_R0_en;
  wire [25:0] mem_23_4_W0_addr;
  wire  mem_23_4_W0_clk;
  wire [7:0] mem_23_4_W0_data;
  wire  mem_23_4_W0_en;
  wire  mem_23_4_W0_mask;
  wire [25:0] mem_23_5_R0_addr;
  wire  mem_23_5_R0_clk;
  wire [7:0] mem_23_5_R0_data;
  wire  mem_23_5_R0_en;
  wire [25:0] mem_23_5_W0_addr;
  wire  mem_23_5_W0_clk;
  wire [7:0] mem_23_5_W0_data;
  wire  mem_23_5_W0_en;
  wire  mem_23_5_W0_mask;
  wire [25:0] mem_23_6_R0_addr;
  wire  mem_23_6_R0_clk;
  wire [7:0] mem_23_6_R0_data;
  wire  mem_23_6_R0_en;
  wire [25:0] mem_23_6_W0_addr;
  wire  mem_23_6_W0_clk;
  wire [7:0] mem_23_6_W0_data;
  wire  mem_23_6_W0_en;
  wire  mem_23_6_W0_mask;
  wire [25:0] mem_23_7_R0_addr;
  wire  mem_23_7_R0_clk;
  wire [7:0] mem_23_7_R0_data;
  wire  mem_23_7_R0_en;
  wire [25:0] mem_23_7_W0_addr;
  wire  mem_23_7_W0_clk;
  wire [7:0] mem_23_7_W0_data;
  wire  mem_23_7_W0_en;
  wire  mem_23_7_W0_mask;
  wire [25:0] mem_24_0_R0_addr;
  wire  mem_24_0_R0_clk;
  wire [7:0] mem_24_0_R0_data;
  wire  mem_24_0_R0_en;
  wire [25:0] mem_24_0_W0_addr;
  wire  mem_24_0_W0_clk;
  wire [7:0] mem_24_0_W0_data;
  wire  mem_24_0_W0_en;
  wire  mem_24_0_W0_mask;
  wire [25:0] mem_24_1_R0_addr;
  wire  mem_24_1_R0_clk;
  wire [7:0] mem_24_1_R0_data;
  wire  mem_24_1_R0_en;
  wire [25:0] mem_24_1_W0_addr;
  wire  mem_24_1_W0_clk;
  wire [7:0] mem_24_1_W0_data;
  wire  mem_24_1_W0_en;
  wire  mem_24_1_W0_mask;
  wire [25:0] mem_24_2_R0_addr;
  wire  mem_24_2_R0_clk;
  wire [7:0] mem_24_2_R0_data;
  wire  mem_24_2_R0_en;
  wire [25:0] mem_24_2_W0_addr;
  wire  mem_24_2_W0_clk;
  wire [7:0] mem_24_2_W0_data;
  wire  mem_24_2_W0_en;
  wire  mem_24_2_W0_mask;
  wire [25:0] mem_24_3_R0_addr;
  wire  mem_24_3_R0_clk;
  wire [7:0] mem_24_3_R0_data;
  wire  mem_24_3_R0_en;
  wire [25:0] mem_24_3_W0_addr;
  wire  mem_24_3_W0_clk;
  wire [7:0] mem_24_3_W0_data;
  wire  mem_24_3_W0_en;
  wire  mem_24_3_W0_mask;
  wire [25:0] mem_24_4_R0_addr;
  wire  mem_24_4_R0_clk;
  wire [7:0] mem_24_4_R0_data;
  wire  mem_24_4_R0_en;
  wire [25:0] mem_24_4_W0_addr;
  wire  mem_24_4_W0_clk;
  wire [7:0] mem_24_4_W0_data;
  wire  mem_24_4_W0_en;
  wire  mem_24_4_W0_mask;
  wire [25:0] mem_24_5_R0_addr;
  wire  mem_24_5_R0_clk;
  wire [7:0] mem_24_5_R0_data;
  wire  mem_24_5_R0_en;
  wire [25:0] mem_24_5_W0_addr;
  wire  mem_24_5_W0_clk;
  wire [7:0] mem_24_5_W0_data;
  wire  mem_24_5_W0_en;
  wire  mem_24_5_W0_mask;
  wire [25:0] mem_24_6_R0_addr;
  wire  mem_24_6_R0_clk;
  wire [7:0] mem_24_6_R0_data;
  wire  mem_24_6_R0_en;
  wire [25:0] mem_24_6_W0_addr;
  wire  mem_24_6_W0_clk;
  wire [7:0] mem_24_6_W0_data;
  wire  mem_24_6_W0_en;
  wire  mem_24_6_W0_mask;
  wire [25:0] mem_24_7_R0_addr;
  wire  mem_24_7_R0_clk;
  wire [7:0] mem_24_7_R0_data;
  wire  mem_24_7_R0_en;
  wire [25:0] mem_24_7_W0_addr;
  wire  mem_24_7_W0_clk;
  wire [7:0] mem_24_7_W0_data;
  wire  mem_24_7_W0_en;
  wire  mem_24_7_W0_mask;
  wire [25:0] mem_25_0_R0_addr;
  wire  mem_25_0_R0_clk;
  wire [7:0] mem_25_0_R0_data;
  wire  mem_25_0_R0_en;
  wire [25:0] mem_25_0_W0_addr;
  wire  mem_25_0_W0_clk;
  wire [7:0] mem_25_0_W0_data;
  wire  mem_25_0_W0_en;
  wire  mem_25_0_W0_mask;
  wire [25:0] mem_25_1_R0_addr;
  wire  mem_25_1_R0_clk;
  wire [7:0] mem_25_1_R0_data;
  wire  mem_25_1_R0_en;
  wire [25:0] mem_25_1_W0_addr;
  wire  mem_25_1_W0_clk;
  wire [7:0] mem_25_1_W0_data;
  wire  mem_25_1_W0_en;
  wire  mem_25_1_W0_mask;
  wire [25:0] mem_25_2_R0_addr;
  wire  mem_25_2_R0_clk;
  wire [7:0] mem_25_2_R0_data;
  wire  mem_25_2_R0_en;
  wire [25:0] mem_25_2_W0_addr;
  wire  mem_25_2_W0_clk;
  wire [7:0] mem_25_2_W0_data;
  wire  mem_25_2_W0_en;
  wire  mem_25_2_W0_mask;
  wire [25:0] mem_25_3_R0_addr;
  wire  mem_25_3_R0_clk;
  wire [7:0] mem_25_3_R0_data;
  wire  mem_25_3_R0_en;
  wire [25:0] mem_25_3_W0_addr;
  wire  mem_25_3_W0_clk;
  wire [7:0] mem_25_3_W0_data;
  wire  mem_25_3_W0_en;
  wire  mem_25_3_W0_mask;
  wire [25:0] mem_25_4_R0_addr;
  wire  mem_25_4_R0_clk;
  wire [7:0] mem_25_4_R0_data;
  wire  mem_25_4_R0_en;
  wire [25:0] mem_25_4_W0_addr;
  wire  mem_25_4_W0_clk;
  wire [7:0] mem_25_4_W0_data;
  wire  mem_25_4_W0_en;
  wire  mem_25_4_W0_mask;
  wire [25:0] mem_25_5_R0_addr;
  wire  mem_25_5_R0_clk;
  wire [7:0] mem_25_5_R0_data;
  wire  mem_25_5_R0_en;
  wire [25:0] mem_25_5_W0_addr;
  wire  mem_25_5_W0_clk;
  wire [7:0] mem_25_5_W0_data;
  wire  mem_25_5_W0_en;
  wire  mem_25_5_W0_mask;
  wire [25:0] mem_25_6_R0_addr;
  wire  mem_25_6_R0_clk;
  wire [7:0] mem_25_6_R0_data;
  wire  mem_25_6_R0_en;
  wire [25:0] mem_25_6_W0_addr;
  wire  mem_25_6_W0_clk;
  wire [7:0] mem_25_6_W0_data;
  wire  mem_25_6_W0_en;
  wire  mem_25_6_W0_mask;
  wire [25:0] mem_25_7_R0_addr;
  wire  mem_25_7_R0_clk;
  wire [7:0] mem_25_7_R0_data;
  wire  mem_25_7_R0_en;
  wire [25:0] mem_25_7_W0_addr;
  wire  mem_25_7_W0_clk;
  wire [7:0] mem_25_7_W0_data;
  wire  mem_25_7_W0_en;
  wire  mem_25_7_W0_mask;
  wire [25:0] mem_26_0_R0_addr;
  wire  mem_26_0_R0_clk;
  wire [7:0] mem_26_0_R0_data;
  wire  mem_26_0_R0_en;
  wire [25:0] mem_26_0_W0_addr;
  wire  mem_26_0_W0_clk;
  wire [7:0] mem_26_0_W0_data;
  wire  mem_26_0_W0_en;
  wire  mem_26_0_W0_mask;
  wire [25:0] mem_26_1_R0_addr;
  wire  mem_26_1_R0_clk;
  wire [7:0] mem_26_1_R0_data;
  wire  mem_26_1_R0_en;
  wire [25:0] mem_26_1_W0_addr;
  wire  mem_26_1_W0_clk;
  wire [7:0] mem_26_1_W0_data;
  wire  mem_26_1_W0_en;
  wire  mem_26_1_W0_mask;
  wire [25:0] mem_26_2_R0_addr;
  wire  mem_26_2_R0_clk;
  wire [7:0] mem_26_2_R0_data;
  wire  mem_26_2_R0_en;
  wire [25:0] mem_26_2_W0_addr;
  wire  mem_26_2_W0_clk;
  wire [7:0] mem_26_2_W0_data;
  wire  mem_26_2_W0_en;
  wire  mem_26_2_W0_mask;
  wire [25:0] mem_26_3_R0_addr;
  wire  mem_26_3_R0_clk;
  wire [7:0] mem_26_3_R0_data;
  wire  mem_26_3_R0_en;
  wire [25:0] mem_26_3_W0_addr;
  wire  mem_26_3_W0_clk;
  wire [7:0] mem_26_3_W0_data;
  wire  mem_26_3_W0_en;
  wire  mem_26_3_W0_mask;
  wire [25:0] mem_26_4_R0_addr;
  wire  mem_26_4_R0_clk;
  wire [7:0] mem_26_4_R0_data;
  wire  mem_26_4_R0_en;
  wire [25:0] mem_26_4_W0_addr;
  wire  mem_26_4_W0_clk;
  wire [7:0] mem_26_4_W0_data;
  wire  mem_26_4_W0_en;
  wire  mem_26_4_W0_mask;
  wire [25:0] mem_26_5_R0_addr;
  wire  mem_26_5_R0_clk;
  wire [7:0] mem_26_5_R0_data;
  wire  mem_26_5_R0_en;
  wire [25:0] mem_26_5_W0_addr;
  wire  mem_26_5_W0_clk;
  wire [7:0] mem_26_5_W0_data;
  wire  mem_26_5_W0_en;
  wire  mem_26_5_W0_mask;
  wire [25:0] mem_26_6_R0_addr;
  wire  mem_26_6_R0_clk;
  wire [7:0] mem_26_6_R0_data;
  wire  mem_26_6_R0_en;
  wire [25:0] mem_26_6_W0_addr;
  wire  mem_26_6_W0_clk;
  wire [7:0] mem_26_6_W0_data;
  wire  mem_26_6_W0_en;
  wire  mem_26_6_W0_mask;
  wire [25:0] mem_26_7_R0_addr;
  wire  mem_26_7_R0_clk;
  wire [7:0] mem_26_7_R0_data;
  wire  mem_26_7_R0_en;
  wire [25:0] mem_26_7_W0_addr;
  wire  mem_26_7_W0_clk;
  wire [7:0] mem_26_7_W0_data;
  wire  mem_26_7_W0_en;
  wire  mem_26_7_W0_mask;
  wire [25:0] mem_27_0_R0_addr;
  wire  mem_27_0_R0_clk;
  wire [7:0] mem_27_0_R0_data;
  wire  mem_27_0_R0_en;
  wire [25:0] mem_27_0_W0_addr;
  wire  mem_27_0_W0_clk;
  wire [7:0] mem_27_0_W0_data;
  wire  mem_27_0_W0_en;
  wire  mem_27_0_W0_mask;
  wire [25:0] mem_27_1_R0_addr;
  wire  mem_27_1_R0_clk;
  wire [7:0] mem_27_1_R0_data;
  wire  mem_27_1_R0_en;
  wire [25:0] mem_27_1_W0_addr;
  wire  mem_27_1_W0_clk;
  wire [7:0] mem_27_1_W0_data;
  wire  mem_27_1_W0_en;
  wire  mem_27_1_W0_mask;
  wire [25:0] mem_27_2_R0_addr;
  wire  mem_27_2_R0_clk;
  wire [7:0] mem_27_2_R0_data;
  wire  mem_27_2_R0_en;
  wire [25:0] mem_27_2_W0_addr;
  wire  mem_27_2_W0_clk;
  wire [7:0] mem_27_2_W0_data;
  wire  mem_27_2_W0_en;
  wire  mem_27_2_W0_mask;
  wire [25:0] mem_27_3_R0_addr;
  wire  mem_27_3_R0_clk;
  wire [7:0] mem_27_3_R0_data;
  wire  mem_27_3_R0_en;
  wire [25:0] mem_27_3_W0_addr;
  wire  mem_27_3_W0_clk;
  wire [7:0] mem_27_3_W0_data;
  wire  mem_27_3_W0_en;
  wire  mem_27_3_W0_mask;
  wire [25:0] mem_27_4_R0_addr;
  wire  mem_27_4_R0_clk;
  wire [7:0] mem_27_4_R0_data;
  wire  mem_27_4_R0_en;
  wire [25:0] mem_27_4_W0_addr;
  wire  mem_27_4_W0_clk;
  wire [7:0] mem_27_4_W0_data;
  wire  mem_27_4_W0_en;
  wire  mem_27_4_W0_mask;
  wire [25:0] mem_27_5_R0_addr;
  wire  mem_27_5_R0_clk;
  wire [7:0] mem_27_5_R0_data;
  wire  mem_27_5_R0_en;
  wire [25:0] mem_27_5_W0_addr;
  wire  mem_27_5_W0_clk;
  wire [7:0] mem_27_5_W0_data;
  wire  mem_27_5_W0_en;
  wire  mem_27_5_W0_mask;
  wire [25:0] mem_27_6_R0_addr;
  wire  mem_27_6_R0_clk;
  wire [7:0] mem_27_6_R0_data;
  wire  mem_27_6_R0_en;
  wire [25:0] mem_27_6_W0_addr;
  wire  mem_27_6_W0_clk;
  wire [7:0] mem_27_6_W0_data;
  wire  mem_27_6_W0_en;
  wire  mem_27_6_W0_mask;
  wire [25:0] mem_27_7_R0_addr;
  wire  mem_27_7_R0_clk;
  wire [7:0] mem_27_7_R0_data;
  wire  mem_27_7_R0_en;
  wire [25:0] mem_27_7_W0_addr;
  wire  mem_27_7_W0_clk;
  wire [7:0] mem_27_7_W0_data;
  wire  mem_27_7_W0_en;
  wire  mem_27_7_W0_mask;
  wire [25:0] mem_28_0_R0_addr;
  wire  mem_28_0_R0_clk;
  wire [7:0] mem_28_0_R0_data;
  wire  mem_28_0_R0_en;
  wire [25:0] mem_28_0_W0_addr;
  wire  mem_28_0_W0_clk;
  wire [7:0] mem_28_0_W0_data;
  wire  mem_28_0_W0_en;
  wire  mem_28_0_W0_mask;
  wire [25:0] mem_28_1_R0_addr;
  wire  mem_28_1_R0_clk;
  wire [7:0] mem_28_1_R0_data;
  wire  mem_28_1_R0_en;
  wire [25:0] mem_28_1_W0_addr;
  wire  mem_28_1_W0_clk;
  wire [7:0] mem_28_1_W0_data;
  wire  mem_28_1_W0_en;
  wire  mem_28_1_W0_mask;
  wire [25:0] mem_28_2_R0_addr;
  wire  mem_28_2_R0_clk;
  wire [7:0] mem_28_2_R0_data;
  wire  mem_28_2_R0_en;
  wire [25:0] mem_28_2_W0_addr;
  wire  mem_28_2_W0_clk;
  wire [7:0] mem_28_2_W0_data;
  wire  mem_28_2_W0_en;
  wire  mem_28_2_W0_mask;
  wire [25:0] mem_28_3_R0_addr;
  wire  mem_28_3_R0_clk;
  wire [7:0] mem_28_3_R0_data;
  wire  mem_28_3_R0_en;
  wire [25:0] mem_28_3_W0_addr;
  wire  mem_28_3_W0_clk;
  wire [7:0] mem_28_3_W0_data;
  wire  mem_28_3_W0_en;
  wire  mem_28_3_W0_mask;
  wire [25:0] mem_28_4_R0_addr;
  wire  mem_28_4_R0_clk;
  wire [7:0] mem_28_4_R0_data;
  wire  mem_28_4_R0_en;
  wire [25:0] mem_28_4_W0_addr;
  wire  mem_28_4_W0_clk;
  wire [7:0] mem_28_4_W0_data;
  wire  mem_28_4_W0_en;
  wire  mem_28_4_W0_mask;
  wire [25:0] mem_28_5_R0_addr;
  wire  mem_28_5_R0_clk;
  wire [7:0] mem_28_5_R0_data;
  wire  mem_28_5_R0_en;
  wire [25:0] mem_28_5_W0_addr;
  wire  mem_28_5_W0_clk;
  wire [7:0] mem_28_5_W0_data;
  wire  mem_28_5_W0_en;
  wire  mem_28_5_W0_mask;
  wire [25:0] mem_28_6_R0_addr;
  wire  mem_28_6_R0_clk;
  wire [7:0] mem_28_6_R0_data;
  wire  mem_28_6_R0_en;
  wire [25:0] mem_28_6_W0_addr;
  wire  mem_28_6_W0_clk;
  wire [7:0] mem_28_6_W0_data;
  wire  mem_28_6_W0_en;
  wire  mem_28_6_W0_mask;
  wire [25:0] mem_28_7_R0_addr;
  wire  mem_28_7_R0_clk;
  wire [7:0] mem_28_7_R0_data;
  wire  mem_28_7_R0_en;
  wire [25:0] mem_28_7_W0_addr;
  wire  mem_28_7_W0_clk;
  wire [7:0] mem_28_7_W0_data;
  wire  mem_28_7_W0_en;
  wire  mem_28_7_W0_mask;
  wire [25:0] mem_29_0_R0_addr;
  wire  mem_29_0_R0_clk;
  wire [7:0] mem_29_0_R0_data;
  wire  mem_29_0_R0_en;
  wire [25:0] mem_29_0_W0_addr;
  wire  mem_29_0_W0_clk;
  wire [7:0] mem_29_0_W0_data;
  wire  mem_29_0_W0_en;
  wire  mem_29_0_W0_mask;
  wire [25:0] mem_29_1_R0_addr;
  wire  mem_29_1_R0_clk;
  wire [7:0] mem_29_1_R0_data;
  wire  mem_29_1_R0_en;
  wire [25:0] mem_29_1_W0_addr;
  wire  mem_29_1_W0_clk;
  wire [7:0] mem_29_1_W0_data;
  wire  mem_29_1_W0_en;
  wire  mem_29_1_W0_mask;
  wire [25:0] mem_29_2_R0_addr;
  wire  mem_29_2_R0_clk;
  wire [7:0] mem_29_2_R0_data;
  wire  mem_29_2_R0_en;
  wire [25:0] mem_29_2_W0_addr;
  wire  mem_29_2_W0_clk;
  wire [7:0] mem_29_2_W0_data;
  wire  mem_29_2_W0_en;
  wire  mem_29_2_W0_mask;
  wire [25:0] mem_29_3_R0_addr;
  wire  mem_29_3_R0_clk;
  wire [7:0] mem_29_3_R0_data;
  wire  mem_29_3_R0_en;
  wire [25:0] mem_29_3_W0_addr;
  wire  mem_29_3_W0_clk;
  wire [7:0] mem_29_3_W0_data;
  wire  mem_29_3_W0_en;
  wire  mem_29_3_W0_mask;
  wire [25:0] mem_29_4_R0_addr;
  wire  mem_29_4_R0_clk;
  wire [7:0] mem_29_4_R0_data;
  wire  mem_29_4_R0_en;
  wire [25:0] mem_29_4_W0_addr;
  wire  mem_29_4_W0_clk;
  wire [7:0] mem_29_4_W0_data;
  wire  mem_29_4_W0_en;
  wire  mem_29_4_W0_mask;
  wire [25:0] mem_29_5_R0_addr;
  wire  mem_29_5_R0_clk;
  wire [7:0] mem_29_5_R0_data;
  wire  mem_29_5_R0_en;
  wire [25:0] mem_29_5_W0_addr;
  wire  mem_29_5_W0_clk;
  wire [7:0] mem_29_5_W0_data;
  wire  mem_29_5_W0_en;
  wire  mem_29_5_W0_mask;
  wire [25:0] mem_29_6_R0_addr;
  wire  mem_29_6_R0_clk;
  wire [7:0] mem_29_6_R0_data;
  wire  mem_29_6_R0_en;
  wire [25:0] mem_29_6_W0_addr;
  wire  mem_29_6_W0_clk;
  wire [7:0] mem_29_6_W0_data;
  wire  mem_29_6_W0_en;
  wire  mem_29_6_W0_mask;
  wire [25:0] mem_29_7_R0_addr;
  wire  mem_29_7_R0_clk;
  wire [7:0] mem_29_7_R0_data;
  wire  mem_29_7_R0_en;
  wire [25:0] mem_29_7_W0_addr;
  wire  mem_29_7_W0_clk;
  wire [7:0] mem_29_7_W0_data;
  wire  mem_29_7_W0_en;
  wire  mem_29_7_W0_mask;
  wire [25:0] mem_30_0_R0_addr;
  wire  mem_30_0_R0_clk;
  wire [7:0] mem_30_0_R0_data;
  wire  mem_30_0_R0_en;
  wire [25:0] mem_30_0_W0_addr;
  wire  mem_30_0_W0_clk;
  wire [7:0] mem_30_0_W0_data;
  wire  mem_30_0_W0_en;
  wire  mem_30_0_W0_mask;
  wire [25:0] mem_30_1_R0_addr;
  wire  mem_30_1_R0_clk;
  wire [7:0] mem_30_1_R0_data;
  wire  mem_30_1_R0_en;
  wire [25:0] mem_30_1_W0_addr;
  wire  mem_30_1_W0_clk;
  wire [7:0] mem_30_1_W0_data;
  wire  mem_30_1_W0_en;
  wire  mem_30_1_W0_mask;
  wire [25:0] mem_30_2_R0_addr;
  wire  mem_30_2_R0_clk;
  wire [7:0] mem_30_2_R0_data;
  wire  mem_30_2_R0_en;
  wire [25:0] mem_30_2_W0_addr;
  wire  mem_30_2_W0_clk;
  wire [7:0] mem_30_2_W0_data;
  wire  mem_30_2_W0_en;
  wire  mem_30_2_W0_mask;
  wire [25:0] mem_30_3_R0_addr;
  wire  mem_30_3_R0_clk;
  wire [7:0] mem_30_3_R0_data;
  wire  mem_30_3_R0_en;
  wire [25:0] mem_30_3_W0_addr;
  wire  mem_30_3_W0_clk;
  wire [7:0] mem_30_3_W0_data;
  wire  mem_30_3_W0_en;
  wire  mem_30_3_W0_mask;
  wire [25:0] mem_30_4_R0_addr;
  wire  mem_30_4_R0_clk;
  wire [7:0] mem_30_4_R0_data;
  wire  mem_30_4_R0_en;
  wire [25:0] mem_30_4_W0_addr;
  wire  mem_30_4_W0_clk;
  wire [7:0] mem_30_4_W0_data;
  wire  mem_30_4_W0_en;
  wire  mem_30_4_W0_mask;
  wire [25:0] mem_30_5_R0_addr;
  wire  mem_30_5_R0_clk;
  wire [7:0] mem_30_5_R0_data;
  wire  mem_30_5_R0_en;
  wire [25:0] mem_30_5_W0_addr;
  wire  mem_30_5_W0_clk;
  wire [7:0] mem_30_5_W0_data;
  wire  mem_30_5_W0_en;
  wire  mem_30_5_W0_mask;
  wire [25:0] mem_30_6_R0_addr;
  wire  mem_30_6_R0_clk;
  wire [7:0] mem_30_6_R0_data;
  wire  mem_30_6_R0_en;
  wire [25:0] mem_30_6_W0_addr;
  wire  mem_30_6_W0_clk;
  wire [7:0] mem_30_6_W0_data;
  wire  mem_30_6_W0_en;
  wire  mem_30_6_W0_mask;
  wire [25:0] mem_30_7_R0_addr;
  wire  mem_30_7_R0_clk;
  wire [7:0] mem_30_7_R0_data;
  wire  mem_30_7_R0_en;
  wire [25:0] mem_30_7_W0_addr;
  wire  mem_30_7_W0_clk;
  wire [7:0] mem_30_7_W0_data;
  wire  mem_30_7_W0_en;
  wire  mem_30_7_W0_mask;
  wire [25:0] mem_31_0_R0_addr;
  wire  mem_31_0_R0_clk;
  wire [7:0] mem_31_0_R0_data;
  wire  mem_31_0_R0_en;
  wire [25:0] mem_31_0_W0_addr;
  wire  mem_31_0_W0_clk;
  wire [7:0] mem_31_0_W0_data;
  wire  mem_31_0_W0_en;
  wire  mem_31_0_W0_mask;
  wire [25:0] mem_31_1_R0_addr;
  wire  mem_31_1_R0_clk;
  wire [7:0] mem_31_1_R0_data;
  wire  mem_31_1_R0_en;
  wire [25:0] mem_31_1_W0_addr;
  wire  mem_31_1_W0_clk;
  wire [7:0] mem_31_1_W0_data;
  wire  mem_31_1_W0_en;
  wire  mem_31_1_W0_mask;
  wire [25:0] mem_31_2_R0_addr;
  wire  mem_31_2_R0_clk;
  wire [7:0] mem_31_2_R0_data;
  wire  mem_31_2_R0_en;
  wire [25:0] mem_31_2_W0_addr;
  wire  mem_31_2_W0_clk;
  wire [7:0] mem_31_2_W0_data;
  wire  mem_31_2_W0_en;
  wire  mem_31_2_W0_mask;
  wire [25:0] mem_31_3_R0_addr;
  wire  mem_31_3_R0_clk;
  wire [7:0] mem_31_3_R0_data;
  wire  mem_31_3_R0_en;
  wire [25:0] mem_31_3_W0_addr;
  wire  mem_31_3_W0_clk;
  wire [7:0] mem_31_3_W0_data;
  wire  mem_31_3_W0_en;
  wire  mem_31_3_W0_mask;
  wire [25:0] mem_31_4_R0_addr;
  wire  mem_31_4_R0_clk;
  wire [7:0] mem_31_4_R0_data;
  wire  mem_31_4_R0_en;
  wire [25:0] mem_31_4_W0_addr;
  wire  mem_31_4_W0_clk;
  wire [7:0] mem_31_4_W0_data;
  wire  mem_31_4_W0_en;
  wire  mem_31_4_W0_mask;
  wire [25:0] mem_31_5_R0_addr;
  wire  mem_31_5_R0_clk;
  wire [7:0] mem_31_5_R0_data;
  wire  mem_31_5_R0_en;
  wire [25:0] mem_31_5_W0_addr;
  wire  mem_31_5_W0_clk;
  wire [7:0] mem_31_5_W0_data;
  wire  mem_31_5_W0_en;
  wire  mem_31_5_W0_mask;
  wire [25:0] mem_31_6_R0_addr;
  wire  mem_31_6_R0_clk;
  wire [7:0] mem_31_6_R0_data;
  wire  mem_31_6_R0_en;
  wire [25:0] mem_31_6_W0_addr;
  wire  mem_31_6_W0_clk;
  wire [7:0] mem_31_6_W0_data;
  wire  mem_31_6_W0_en;
  wire  mem_31_6_W0_mask;
  wire [25:0] mem_31_7_R0_addr;
  wire  mem_31_7_R0_clk;
  wire [7:0] mem_31_7_R0_data;
  wire  mem_31_7_R0_en;
  wire [25:0] mem_31_7_W0_addr;
  wire  mem_31_7_W0_clk;
  wire [7:0] mem_31_7_W0_data;
  wire  mem_31_7_W0_en;
  wire  mem_31_7_W0_mask;
  wire [25:0] mem_32_0_R0_addr;
  wire  mem_32_0_R0_clk;
  wire [7:0] mem_32_0_R0_data;
  wire  mem_32_0_R0_en;
  wire [25:0] mem_32_0_W0_addr;
  wire  mem_32_0_W0_clk;
  wire [7:0] mem_32_0_W0_data;
  wire  mem_32_0_W0_en;
  wire  mem_32_0_W0_mask;
  wire [25:0] mem_32_1_R0_addr;
  wire  mem_32_1_R0_clk;
  wire [7:0] mem_32_1_R0_data;
  wire  mem_32_1_R0_en;
  wire [25:0] mem_32_1_W0_addr;
  wire  mem_32_1_W0_clk;
  wire [7:0] mem_32_1_W0_data;
  wire  mem_32_1_W0_en;
  wire  mem_32_1_W0_mask;
  wire [25:0] mem_32_2_R0_addr;
  wire  mem_32_2_R0_clk;
  wire [7:0] mem_32_2_R0_data;
  wire  mem_32_2_R0_en;
  wire [25:0] mem_32_2_W0_addr;
  wire  mem_32_2_W0_clk;
  wire [7:0] mem_32_2_W0_data;
  wire  mem_32_2_W0_en;
  wire  mem_32_2_W0_mask;
  wire [25:0] mem_32_3_R0_addr;
  wire  mem_32_3_R0_clk;
  wire [7:0] mem_32_3_R0_data;
  wire  mem_32_3_R0_en;
  wire [25:0] mem_32_3_W0_addr;
  wire  mem_32_3_W0_clk;
  wire [7:0] mem_32_3_W0_data;
  wire  mem_32_3_W0_en;
  wire  mem_32_3_W0_mask;
  wire [25:0] mem_32_4_R0_addr;
  wire  mem_32_4_R0_clk;
  wire [7:0] mem_32_4_R0_data;
  wire  mem_32_4_R0_en;
  wire [25:0] mem_32_4_W0_addr;
  wire  mem_32_4_W0_clk;
  wire [7:0] mem_32_4_W0_data;
  wire  mem_32_4_W0_en;
  wire  mem_32_4_W0_mask;
  wire [25:0] mem_32_5_R0_addr;
  wire  mem_32_5_R0_clk;
  wire [7:0] mem_32_5_R0_data;
  wire  mem_32_5_R0_en;
  wire [25:0] mem_32_5_W0_addr;
  wire  mem_32_5_W0_clk;
  wire [7:0] mem_32_5_W0_data;
  wire  mem_32_5_W0_en;
  wire  mem_32_5_W0_mask;
  wire [25:0] mem_32_6_R0_addr;
  wire  mem_32_6_R0_clk;
  wire [7:0] mem_32_6_R0_data;
  wire  mem_32_6_R0_en;
  wire [25:0] mem_32_6_W0_addr;
  wire  mem_32_6_W0_clk;
  wire [7:0] mem_32_6_W0_data;
  wire  mem_32_6_W0_en;
  wire  mem_32_6_W0_mask;
  wire [25:0] mem_32_7_R0_addr;
  wire  mem_32_7_R0_clk;
  wire [7:0] mem_32_7_R0_data;
  wire  mem_32_7_R0_en;
  wire [25:0] mem_32_7_W0_addr;
  wire  mem_32_7_W0_clk;
  wire [7:0] mem_32_7_W0_data;
  wire  mem_32_7_W0_en;
  wire  mem_32_7_W0_mask;
  wire [25:0] mem_33_0_R0_addr;
  wire  mem_33_0_R0_clk;
  wire [7:0] mem_33_0_R0_data;
  wire  mem_33_0_R0_en;
  wire [25:0] mem_33_0_W0_addr;
  wire  mem_33_0_W0_clk;
  wire [7:0] mem_33_0_W0_data;
  wire  mem_33_0_W0_en;
  wire  mem_33_0_W0_mask;
  wire [25:0] mem_33_1_R0_addr;
  wire  mem_33_1_R0_clk;
  wire [7:0] mem_33_1_R0_data;
  wire  mem_33_1_R0_en;
  wire [25:0] mem_33_1_W0_addr;
  wire  mem_33_1_W0_clk;
  wire [7:0] mem_33_1_W0_data;
  wire  mem_33_1_W0_en;
  wire  mem_33_1_W0_mask;
  wire [25:0] mem_33_2_R0_addr;
  wire  mem_33_2_R0_clk;
  wire [7:0] mem_33_2_R0_data;
  wire  mem_33_2_R0_en;
  wire [25:0] mem_33_2_W0_addr;
  wire  mem_33_2_W0_clk;
  wire [7:0] mem_33_2_W0_data;
  wire  mem_33_2_W0_en;
  wire  mem_33_2_W0_mask;
  wire [25:0] mem_33_3_R0_addr;
  wire  mem_33_3_R0_clk;
  wire [7:0] mem_33_3_R0_data;
  wire  mem_33_3_R0_en;
  wire [25:0] mem_33_3_W0_addr;
  wire  mem_33_3_W0_clk;
  wire [7:0] mem_33_3_W0_data;
  wire  mem_33_3_W0_en;
  wire  mem_33_3_W0_mask;
  wire [25:0] mem_33_4_R0_addr;
  wire  mem_33_4_R0_clk;
  wire [7:0] mem_33_4_R0_data;
  wire  mem_33_4_R0_en;
  wire [25:0] mem_33_4_W0_addr;
  wire  mem_33_4_W0_clk;
  wire [7:0] mem_33_4_W0_data;
  wire  mem_33_4_W0_en;
  wire  mem_33_4_W0_mask;
  wire [25:0] mem_33_5_R0_addr;
  wire  mem_33_5_R0_clk;
  wire [7:0] mem_33_5_R0_data;
  wire  mem_33_5_R0_en;
  wire [25:0] mem_33_5_W0_addr;
  wire  mem_33_5_W0_clk;
  wire [7:0] mem_33_5_W0_data;
  wire  mem_33_5_W0_en;
  wire  mem_33_5_W0_mask;
  wire [25:0] mem_33_6_R0_addr;
  wire  mem_33_6_R0_clk;
  wire [7:0] mem_33_6_R0_data;
  wire  mem_33_6_R0_en;
  wire [25:0] mem_33_6_W0_addr;
  wire  mem_33_6_W0_clk;
  wire [7:0] mem_33_6_W0_data;
  wire  mem_33_6_W0_en;
  wire  mem_33_6_W0_mask;
  wire [25:0] mem_33_7_R0_addr;
  wire  mem_33_7_R0_clk;
  wire [7:0] mem_33_7_R0_data;
  wire  mem_33_7_R0_en;
  wire [25:0] mem_33_7_W0_addr;
  wire  mem_33_7_W0_clk;
  wire [7:0] mem_33_7_W0_data;
  wire  mem_33_7_W0_en;
  wire  mem_33_7_W0_mask;
  wire [25:0] mem_34_0_R0_addr;
  wire  mem_34_0_R0_clk;
  wire [7:0] mem_34_0_R0_data;
  wire  mem_34_0_R0_en;
  wire [25:0] mem_34_0_W0_addr;
  wire  mem_34_0_W0_clk;
  wire [7:0] mem_34_0_W0_data;
  wire  mem_34_0_W0_en;
  wire  mem_34_0_W0_mask;
  wire [25:0] mem_34_1_R0_addr;
  wire  mem_34_1_R0_clk;
  wire [7:0] mem_34_1_R0_data;
  wire  mem_34_1_R0_en;
  wire [25:0] mem_34_1_W0_addr;
  wire  mem_34_1_W0_clk;
  wire [7:0] mem_34_1_W0_data;
  wire  mem_34_1_W0_en;
  wire  mem_34_1_W0_mask;
  wire [25:0] mem_34_2_R0_addr;
  wire  mem_34_2_R0_clk;
  wire [7:0] mem_34_2_R0_data;
  wire  mem_34_2_R0_en;
  wire [25:0] mem_34_2_W0_addr;
  wire  mem_34_2_W0_clk;
  wire [7:0] mem_34_2_W0_data;
  wire  mem_34_2_W0_en;
  wire  mem_34_2_W0_mask;
  wire [25:0] mem_34_3_R0_addr;
  wire  mem_34_3_R0_clk;
  wire [7:0] mem_34_3_R0_data;
  wire  mem_34_3_R0_en;
  wire [25:0] mem_34_3_W0_addr;
  wire  mem_34_3_W0_clk;
  wire [7:0] mem_34_3_W0_data;
  wire  mem_34_3_W0_en;
  wire  mem_34_3_W0_mask;
  wire [25:0] mem_34_4_R0_addr;
  wire  mem_34_4_R0_clk;
  wire [7:0] mem_34_4_R0_data;
  wire  mem_34_4_R0_en;
  wire [25:0] mem_34_4_W0_addr;
  wire  mem_34_4_W0_clk;
  wire [7:0] mem_34_4_W0_data;
  wire  mem_34_4_W0_en;
  wire  mem_34_4_W0_mask;
  wire [25:0] mem_34_5_R0_addr;
  wire  mem_34_5_R0_clk;
  wire [7:0] mem_34_5_R0_data;
  wire  mem_34_5_R0_en;
  wire [25:0] mem_34_5_W0_addr;
  wire  mem_34_5_W0_clk;
  wire [7:0] mem_34_5_W0_data;
  wire  mem_34_5_W0_en;
  wire  mem_34_5_W0_mask;
  wire [25:0] mem_34_6_R0_addr;
  wire  mem_34_6_R0_clk;
  wire [7:0] mem_34_6_R0_data;
  wire  mem_34_6_R0_en;
  wire [25:0] mem_34_6_W0_addr;
  wire  mem_34_6_W0_clk;
  wire [7:0] mem_34_6_W0_data;
  wire  mem_34_6_W0_en;
  wire  mem_34_6_W0_mask;
  wire [25:0] mem_34_7_R0_addr;
  wire  mem_34_7_R0_clk;
  wire [7:0] mem_34_7_R0_data;
  wire  mem_34_7_R0_en;
  wire [25:0] mem_34_7_W0_addr;
  wire  mem_34_7_W0_clk;
  wire [7:0] mem_34_7_W0_data;
  wire  mem_34_7_W0_en;
  wire  mem_34_7_W0_mask;
  wire [25:0] mem_35_0_R0_addr;
  wire  mem_35_0_R0_clk;
  wire [7:0] mem_35_0_R0_data;
  wire  mem_35_0_R0_en;
  wire [25:0] mem_35_0_W0_addr;
  wire  mem_35_0_W0_clk;
  wire [7:0] mem_35_0_W0_data;
  wire  mem_35_0_W0_en;
  wire  mem_35_0_W0_mask;
  wire [25:0] mem_35_1_R0_addr;
  wire  mem_35_1_R0_clk;
  wire [7:0] mem_35_1_R0_data;
  wire  mem_35_1_R0_en;
  wire [25:0] mem_35_1_W0_addr;
  wire  mem_35_1_W0_clk;
  wire [7:0] mem_35_1_W0_data;
  wire  mem_35_1_W0_en;
  wire  mem_35_1_W0_mask;
  wire [25:0] mem_35_2_R0_addr;
  wire  mem_35_2_R0_clk;
  wire [7:0] mem_35_2_R0_data;
  wire  mem_35_2_R0_en;
  wire [25:0] mem_35_2_W0_addr;
  wire  mem_35_2_W0_clk;
  wire [7:0] mem_35_2_W0_data;
  wire  mem_35_2_W0_en;
  wire  mem_35_2_W0_mask;
  wire [25:0] mem_35_3_R0_addr;
  wire  mem_35_3_R0_clk;
  wire [7:0] mem_35_3_R0_data;
  wire  mem_35_3_R0_en;
  wire [25:0] mem_35_3_W0_addr;
  wire  mem_35_3_W0_clk;
  wire [7:0] mem_35_3_W0_data;
  wire  mem_35_3_W0_en;
  wire  mem_35_3_W0_mask;
  wire [25:0] mem_35_4_R0_addr;
  wire  mem_35_4_R0_clk;
  wire [7:0] mem_35_4_R0_data;
  wire  mem_35_4_R0_en;
  wire [25:0] mem_35_4_W0_addr;
  wire  mem_35_4_W0_clk;
  wire [7:0] mem_35_4_W0_data;
  wire  mem_35_4_W0_en;
  wire  mem_35_4_W0_mask;
  wire [25:0] mem_35_5_R0_addr;
  wire  mem_35_5_R0_clk;
  wire [7:0] mem_35_5_R0_data;
  wire  mem_35_5_R0_en;
  wire [25:0] mem_35_5_W0_addr;
  wire  mem_35_5_W0_clk;
  wire [7:0] mem_35_5_W0_data;
  wire  mem_35_5_W0_en;
  wire  mem_35_5_W0_mask;
  wire [25:0] mem_35_6_R0_addr;
  wire  mem_35_6_R0_clk;
  wire [7:0] mem_35_6_R0_data;
  wire  mem_35_6_R0_en;
  wire [25:0] mem_35_6_W0_addr;
  wire  mem_35_6_W0_clk;
  wire [7:0] mem_35_6_W0_data;
  wire  mem_35_6_W0_en;
  wire  mem_35_6_W0_mask;
  wire [25:0] mem_35_7_R0_addr;
  wire  mem_35_7_R0_clk;
  wire [7:0] mem_35_7_R0_data;
  wire  mem_35_7_R0_en;
  wire [25:0] mem_35_7_W0_addr;
  wire  mem_35_7_W0_clk;
  wire [7:0] mem_35_7_W0_data;
  wire  mem_35_7_W0_en;
  wire  mem_35_7_W0_mask;
  wire [25:0] mem_36_0_R0_addr;
  wire  mem_36_0_R0_clk;
  wire [7:0] mem_36_0_R0_data;
  wire  mem_36_0_R0_en;
  wire [25:0] mem_36_0_W0_addr;
  wire  mem_36_0_W0_clk;
  wire [7:0] mem_36_0_W0_data;
  wire  mem_36_0_W0_en;
  wire  mem_36_0_W0_mask;
  wire [25:0] mem_36_1_R0_addr;
  wire  mem_36_1_R0_clk;
  wire [7:0] mem_36_1_R0_data;
  wire  mem_36_1_R0_en;
  wire [25:0] mem_36_1_W0_addr;
  wire  mem_36_1_W0_clk;
  wire [7:0] mem_36_1_W0_data;
  wire  mem_36_1_W0_en;
  wire  mem_36_1_W0_mask;
  wire [25:0] mem_36_2_R0_addr;
  wire  mem_36_2_R0_clk;
  wire [7:0] mem_36_2_R0_data;
  wire  mem_36_2_R0_en;
  wire [25:0] mem_36_2_W0_addr;
  wire  mem_36_2_W0_clk;
  wire [7:0] mem_36_2_W0_data;
  wire  mem_36_2_W0_en;
  wire  mem_36_2_W0_mask;
  wire [25:0] mem_36_3_R0_addr;
  wire  mem_36_3_R0_clk;
  wire [7:0] mem_36_3_R0_data;
  wire  mem_36_3_R0_en;
  wire [25:0] mem_36_3_W0_addr;
  wire  mem_36_3_W0_clk;
  wire [7:0] mem_36_3_W0_data;
  wire  mem_36_3_W0_en;
  wire  mem_36_3_W0_mask;
  wire [25:0] mem_36_4_R0_addr;
  wire  mem_36_4_R0_clk;
  wire [7:0] mem_36_4_R0_data;
  wire  mem_36_4_R0_en;
  wire [25:0] mem_36_4_W0_addr;
  wire  mem_36_4_W0_clk;
  wire [7:0] mem_36_4_W0_data;
  wire  mem_36_4_W0_en;
  wire  mem_36_4_W0_mask;
  wire [25:0] mem_36_5_R0_addr;
  wire  mem_36_5_R0_clk;
  wire [7:0] mem_36_5_R0_data;
  wire  mem_36_5_R0_en;
  wire [25:0] mem_36_5_W0_addr;
  wire  mem_36_5_W0_clk;
  wire [7:0] mem_36_5_W0_data;
  wire  mem_36_5_W0_en;
  wire  mem_36_5_W0_mask;
  wire [25:0] mem_36_6_R0_addr;
  wire  mem_36_6_R0_clk;
  wire [7:0] mem_36_6_R0_data;
  wire  mem_36_6_R0_en;
  wire [25:0] mem_36_6_W0_addr;
  wire  mem_36_6_W0_clk;
  wire [7:0] mem_36_6_W0_data;
  wire  mem_36_6_W0_en;
  wire  mem_36_6_W0_mask;
  wire [25:0] mem_36_7_R0_addr;
  wire  mem_36_7_R0_clk;
  wire [7:0] mem_36_7_R0_data;
  wire  mem_36_7_R0_en;
  wire [25:0] mem_36_7_W0_addr;
  wire  mem_36_7_W0_clk;
  wire [7:0] mem_36_7_W0_data;
  wire  mem_36_7_W0_en;
  wire  mem_36_7_W0_mask;
  wire [25:0] mem_37_0_R0_addr;
  wire  mem_37_0_R0_clk;
  wire [7:0] mem_37_0_R0_data;
  wire  mem_37_0_R0_en;
  wire [25:0] mem_37_0_W0_addr;
  wire  mem_37_0_W0_clk;
  wire [7:0] mem_37_0_W0_data;
  wire  mem_37_0_W0_en;
  wire  mem_37_0_W0_mask;
  wire [25:0] mem_37_1_R0_addr;
  wire  mem_37_1_R0_clk;
  wire [7:0] mem_37_1_R0_data;
  wire  mem_37_1_R0_en;
  wire [25:0] mem_37_1_W0_addr;
  wire  mem_37_1_W0_clk;
  wire [7:0] mem_37_1_W0_data;
  wire  mem_37_1_W0_en;
  wire  mem_37_1_W0_mask;
  wire [25:0] mem_37_2_R0_addr;
  wire  mem_37_2_R0_clk;
  wire [7:0] mem_37_2_R0_data;
  wire  mem_37_2_R0_en;
  wire [25:0] mem_37_2_W0_addr;
  wire  mem_37_2_W0_clk;
  wire [7:0] mem_37_2_W0_data;
  wire  mem_37_2_W0_en;
  wire  mem_37_2_W0_mask;
  wire [25:0] mem_37_3_R0_addr;
  wire  mem_37_3_R0_clk;
  wire [7:0] mem_37_3_R0_data;
  wire  mem_37_3_R0_en;
  wire [25:0] mem_37_3_W0_addr;
  wire  mem_37_3_W0_clk;
  wire [7:0] mem_37_3_W0_data;
  wire  mem_37_3_W0_en;
  wire  mem_37_3_W0_mask;
  wire [25:0] mem_37_4_R0_addr;
  wire  mem_37_4_R0_clk;
  wire [7:0] mem_37_4_R0_data;
  wire  mem_37_4_R0_en;
  wire [25:0] mem_37_4_W0_addr;
  wire  mem_37_4_W0_clk;
  wire [7:0] mem_37_4_W0_data;
  wire  mem_37_4_W0_en;
  wire  mem_37_4_W0_mask;
  wire [25:0] mem_37_5_R0_addr;
  wire  mem_37_5_R0_clk;
  wire [7:0] mem_37_5_R0_data;
  wire  mem_37_5_R0_en;
  wire [25:0] mem_37_5_W0_addr;
  wire  mem_37_5_W0_clk;
  wire [7:0] mem_37_5_W0_data;
  wire  mem_37_5_W0_en;
  wire  mem_37_5_W0_mask;
  wire [25:0] mem_37_6_R0_addr;
  wire  mem_37_6_R0_clk;
  wire [7:0] mem_37_6_R0_data;
  wire  mem_37_6_R0_en;
  wire [25:0] mem_37_6_W0_addr;
  wire  mem_37_6_W0_clk;
  wire [7:0] mem_37_6_W0_data;
  wire  mem_37_6_W0_en;
  wire  mem_37_6_W0_mask;
  wire [25:0] mem_37_7_R0_addr;
  wire  mem_37_7_R0_clk;
  wire [7:0] mem_37_7_R0_data;
  wire  mem_37_7_R0_en;
  wire [25:0] mem_37_7_W0_addr;
  wire  mem_37_7_W0_clk;
  wire [7:0] mem_37_7_W0_data;
  wire  mem_37_7_W0_en;
  wire  mem_37_7_W0_mask;
  wire [25:0] mem_38_0_R0_addr;
  wire  mem_38_0_R0_clk;
  wire [7:0] mem_38_0_R0_data;
  wire  mem_38_0_R0_en;
  wire [25:0] mem_38_0_W0_addr;
  wire  mem_38_0_W0_clk;
  wire [7:0] mem_38_0_W0_data;
  wire  mem_38_0_W0_en;
  wire  mem_38_0_W0_mask;
  wire [25:0] mem_38_1_R0_addr;
  wire  mem_38_1_R0_clk;
  wire [7:0] mem_38_1_R0_data;
  wire  mem_38_1_R0_en;
  wire [25:0] mem_38_1_W0_addr;
  wire  mem_38_1_W0_clk;
  wire [7:0] mem_38_1_W0_data;
  wire  mem_38_1_W0_en;
  wire  mem_38_1_W0_mask;
  wire [25:0] mem_38_2_R0_addr;
  wire  mem_38_2_R0_clk;
  wire [7:0] mem_38_2_R0_data;
  wire  mem_38_2_R0_en;
  wire [25:0] mem_38_2_W0_addr;
  wire  mem_38_2_W0_clk;
  wire [7:0] mem_38_2_W0_data;
  wire  mem_38_2_W0_en;
  wire  mem_38_2_W0_mask;
  wire [25:0] mem_38_3_R0_addr;
  wire  mem_38_3_R0_clk;
  wire [7:0] mem_38_3_R0_data;
  wire  mem_38_3_R0_en;
  wire [25:0] mem_38_3_W0_addr;
  wire  mem_38_3_W0_clk;
  wire [7:0] mem_38_3_W0_data;
  wire  mem_38_3_W0_en;
  wire  mem_38_3_W0_mask;
  wire [25:0] mem_38_4_R0_addr;
  wire  mem_38_4_R0_clk;
  wire [7:0] mem_38_4_R0_data;
  wire  mem_38_4_R0_en;
  wire [25:0] mem_38_4_W0_addr;
  wire  mem_38_4_W0_clk;
  wire [7:0] mem_38_4_W0_data;
  wire  mem_38_4_W0_en;
  wire  mem_38_4_W0_mask;
  wire [25:0] mem_38_5_R0_addr;
  wire  mem_38_5_R0_clk;
  wire [7:0] mem_38_5_R0_data;
  wire  mem_38_5_R0_en;
  wire [25:0] mem_38_5_W0_addr;
  wire  mem_38_5_W0_clk;
  wire [7:0] mem_38_5_W0_data;
  wire  mem_38_5_W0_en;
  wire  mem_38_5_W0_mask;
  wire [25:0] mem_38_6_R0_addr;
  wire  mem_38_6_R0_clk;
  wire [7:0] mem_38_6_R0_data;
  wire  mem_38_6_R0_en;
  wire [25:0] mem_38_6_W0_addr;
  wire  mem_38_6_W0_clk;
  wire [7:0] mem_38_6_W0_data;
  wire  mem_38_6_W0_en;
  wire  mem_38_6_W0_mask;
  wire [25:0] mem_38_7_R0_addr;
  wire  mem_38_7_R0_clk;
  wire [7:0] mem_38_7_R0_data;
  wire  mem_38_7_R0_en;
  wire [25:0] mem_38_7_W0_addr;
  wire  mem_38_7_W0_clk;
  wire [7:0] mem_38_7_W0_data;
  wire  mem_38_7_W0_en;
  wire  mem_38_7_W0_mask;
  wire [25:0] mem_39_0_R0_addr;
  wire  mem_39_0_R0_clk;
  wire [7:0] mem_39_0_R0_data;
  wire  mem_39_0_R0_en;
  wire [25:0] mem_39_0_W0_addr;
  wire  mem_39_0_W0_clk;
  wire [7:0] mem_39_0_W0_data;
  wire  mem_39_0_W0_en;
  wire  mem_39_0_W0_mask;
  wire [25:0] mem_39_1_R0_addr;
  wire  mem_39_1_R0_clk;
  wire [7:0] mem_39_1_R0_data;
  wire  mem_39_1_R0_en;
  wire [25:0] mem_39_1_W0_addr;
  wire  mem_39_1_W0_clk;
  wire [7:0] mem_39_1_W0_data;
  wire  mem_39_1_W0_en;
  wire  mem_39_1_W0_mask;
  wire [25:0] mem_39_2_R0_addr;
  wire  mem_39_2_R0_clk;
  wire [7:0] mem_39_2_R0_data;
  wire  mem_39_2_R0_en;
  wire [25:0] mem_39_2_W0_addr;
  wire  mem_39_2_W0_clk;
  wire [7:0] mem_39_2_W0_data;
  wire  mem_39_2_W0_en;
  wire  mem_39_2_W0_mask;
  wire [25:0] mem_39_3_R0_addr;
  wire  mem_39_3_R0_clk;
  wire [7:0] mem_39_3_R0_data;
  wire  mem_39_3_R0_en;
  wire [25:0] mem_39_3_W0_addr;
  wire  mem_39_3_W0_clk;
  wire [7:0] mem_39_3_W0_data;
  wire  mem_39_3_W0_en;
  wire  mem_39_3_W0_mask;
  wire [25:0] mem_39_4_R0_addr;
  wire  mem_39_4_R0_clk;
  wire [7:0] mem_39_4_R0_data;
  wire  mem_39_4_R0_en;
  wire [25:0] mem_39_4_W0_addr;
  wire  mem_39_4_W0_clk;
  wire [7:0] mem_39_4_W0_data;
  wire  mem_39_4_W0_en;
  wire  mem_39_4_W0_mask;
  wire [25:0] mem_39_5_R0_addr;
  wire  mem_39_5_R0_clk;
  wire [7:0] mem_39_5_R0_data;
  wire  mem_39_5_R0_en;
  wire [25:0] mem_39_5_W0_addr;
  wire  mem_39_5_W0_clk;
  wire [7:0] mem_39_5_W0_data;
  wire  mem_39_5_W0_en;
  wire  mem_39_5_W0_mask;
  wire [25:0] mem_39_6_R0_addr;
  wire  mem_39_6_R0_clk;
  wire [7:0] mem_39_6_R0_data;
  wire  mem_39_6_R0_en;
  wire [25:0] mem_39_6_W0_addr;
  wire  mem_39_6_W0_clk;
  wire [7:0] mem_39_6_W0_data;
  wire  mem_39_6_W0_en;
  wire  mem_39_6_W0_mask;
  wire [25:0] mem_39_7_R0_addr;
  wire  mem_39_7_R0_clk;
  wire [7:0] mem_39_7_R0_data;
  wire  mem_39_7_R0_en;
  wire [25:0] mem_39_7_W0_addr;
  wire  mem_39_7_W0_clk;
  wire [7:0] mem_39_7_W0_data;
  wire  mem_39_7_W0_en;
  wire  mem_39_7_W0_mask;
  wire [25:0] mem_40_0_R0_addr;
  wire  mem_40_0_R0_clk;
  wire [7:0] mem_40_0_R0_data;
  wire  mem_40_0_R0_en;
  wire [25:0] mem_40_0_W0_addr;
  wire  mem_40_0_W0_clk;
  wire [7:0] mem_40_0_W0_data;
  wire  mem_40_0_W0_en;
  wire  mem_40_0_W0_mask;
  wire [25:0] mem_40_1_R0_addr;
  wire  mem_40_1_R0_clk;
  wire [7:0] mem_40_1_R0_data;
  wire  mem_40_1_R0_en;
  wire [25:0] mem_40_1_W0_addr;
  wire  mem_40_1_W0_clk;
  wire [7:0] mem_40_1_W0_data;
  wire  mem_40_1_W0_en;
  wire  mem_40_1_W0_mask;
  wire [25:0] mem_40_2_R0_addr;
  wire  mem_40_2_R0_clk;
  wire [7:0] mem_40_2_R0_data;
  wire  mem_40_2_R0_en;
  wire [25:0] mem_40_2_W0_addr;
  wire  mem_40_2_W0_clk;
  wire [7:0] mem_40_2_W0_data;
  wire  mem_40_2_W0_en;
  wire  mem_40_2_W0_mask;
  wire [25:0] mem_40_3_R0_addr;
  wire  mem_40_3_R0_clk;
  wire [7:0] mem_40_3_R0_data;
  wire  mem_40_3_R0_en;
  wire [25:0] mem_40_3_W0_addr;
  wire  mem_40_3_W0_clk;
  wire [7:0] mem_40_3_W0_data;
  wire  mem_40_3_W0_en;
  wire  mem_40_3_W0_mask;
  wire [25:0] mem_40_4_R0_addr;
  wire  mem_40_4_R0_clk;
  wire [7:0] mem_40_4_R0_data;
  wire  mem_40_4_R0_en;
  wire [25:0] mem_40_4_W0_addr;
  wire  mem_40_4_W0_clk;
  wire [7:0] mem_40_4_W0_data;
  wire  mem_40_4_W0_en;
  wire  mem_40_4_W0_mask;
  wire [25:0] mem_40_5_R0_addr;
  wire  mem_40_5_R0_clk;
  wire [7:0] mem_40_5_R0_data;
  wire  mem_40_5_R0_en;
  wire [25:0] mem_40_5_W0_addr;
  wire  mem_40_5_W0_clk;
  wire [7:0] mem_40_5_W0_data;
  wire  mem_40_5_W0_en;
  wire  mem_40_5_W0_mask;
  wire [25:0] mem_40_6_R0_addr;
  wire  mem_40_6_R0_clk;
  wire [7:0] mem_40_6_R0_data;
  wire  mem_40_6_R0_en;
  wire [25:0] mem_40_6_W0_addr;
  wire  mem_40_6_W0_clk;
  wire [7:0] mem_40_6_W0_data;
  wire  mem_40_6_W0_en;
  wire  mem_40_6_W0_mask;
  wire [25:0] mem_40_7_R0_addr;
  wire  mem_40_7_R0_clk;
  wire [7:0] mem_40_7_R0_data;
  wire  mem_40_7_R0_en;
  wire [25:0] mem_40_7_W0_addr;
  wire  mem_40_7_W0_clk;
  wire [7:0] mem_40_7_W0_data;
  wire  mem_40_7_W0_en;
  wire  mem_40_7_W0_mask;
  wire [25:0] mem_41_0_R0_addr;
  wire  mem_41_0_R0_clk;
  wire [7:0] mem_41_0_R0_data;
  wire  mem_41_0_R0_en;
  wire [25:0] mem_41_0_W0_addr;
  wire  mem_41_0_W0_clk;
  wire [7:0] mem_41_0_W0_data;
  wire  mem_41_0_W0_en;
  wire  mem_41_0_W0_mask;
  wire [25:0] mem_41_1_R0_addr;
  wire  mem_41_1_R0_clk;
  wire [7:0] mem_41_1_R0_data;
  wire  mem_41_1_R0_en;
  wire [25:0] mem_41_1_W0_addr;
  wire  mem_41_1_W0_clk;
  wire [7:0] mem_41_1_W0_data;
  wire  mem_41_1_W0_en;
  wire  mem_41_1_W0_mask;
  wire [25:0] mem_41_2_R0_addr;
  wire  mem_41_2_R0_clk;
  wire [7:0] mem_41_2_R0_data;
  wire  mem_41_2_R0_en;
  wire [25:0] mem_41_2_W0_addr;
  wire  mem_41_2_W0_clk;
  wire [7:0] mem_41_2_W0_data;
  wire  mem_41_2_W0_en;
  wire  mem_41_2_W0_mask;
  wire [25:0] mem_41_3_R0_addr;
  wire  mem_41_3_R0_clk;
  wire [7:0] mem_41_3_R0_data;
  wire  mem_41_3_R0_en;
  wire [25:0] mem_41_3_W0_addr;
  wire  mem_41_3_W0_clk;
  wire [7:0] mem_41_3_W0_data;
  wire  mem_41_3_W0_en;
  wire  mem_41_3_W0_mask;
  wire [25:0] mem_41_4_R0_addr;
  wire  mem_41_4_R0_clk;
  wire [7:0] mem_41_4_R0_data;
  wire  mem_41_4_R0_en;
  wire [25:0] mem_41_4_W0_addr;
  wire  mem_41_4_W0_clk;
  wire [7:0] mem_41_4_W0_data;
  wire  mem_41_4_W0_en;
  wire  mem_41_4_W0_mask;
  wire [25:0] mem_41_5_R0_addr;
  wire  mem_41_5_R0_clk;
  wire [7:0] mem_41_5_R0_data;
  wire  mem_41_5_R0_en;
  wire [25:0] mem_41_5_W0_addr;
  wire  mem_41_5_W0_clk;
  wire [7:0] mem_41_5_W0_data;
  wire  mem_41_5_W0_en;
  wire  mem_41_5_W0_mask;
  wire [25:0] mem_41_6_R0_addr;
  wire  mem_41_6_R0_clk;
  wire [7:0] mem_41_6_R0_data;
  wire  mem_41_6_R0_en;
  wire [25:0] mem_41_6_W0_addr;
  wire  mem_41_6_W0_clk;
  wire [7:0] mem_41_6_W0_data;
  wire  mem_41_6_W0_en;
  wire  mem_41_6_W0_mask;
  wire [25:0] mem_41_7_R0_addr;
  wire  mem_41_7_R0_clk;
  wire [7:0] mem_41_7_R0_data;
  wire  mem_41_7_R0_en;
  wire [25:0] mem_41_7_W0_addr;
  wire  mem_41_7_W0_clk;
  wire [7:0] mem_41_7_W0_data;
  wire  mem_41_7_W0_en;
  wire  mem_41_7_W0_mask;
  wire [25:0] mem_42_0_R0_addr;
  wire  mem_42_0_R0_clk;
  wire [7:0] mem_42_0_R0_data;
  wire  mem_42_0_R0_en;
  wire [25:0] mem_42_0_W0_addr;
  wire  mem_42_0_W0_clk;
  wire [7:0] mem_42_0_W0_data;
  wire  mem_42_0_W0_en;
  wire  mem_42_0_W0_mask;
  wire [25:0] mem_42_1_R0_addr;
  wire  mem_42_1_R0_clk;
  wire [7:0] mem_42_1_R0_data;
  wire  mem_42_1_R0_en;
  wire [25:0] mem_42_1_W0_addr;
  wire  mem_42_1_W0_clk;
  wire [7:0] mem_42_1_W0_data;
  wire  mem_42_1_W0_en;
  wire  mem_42_1_W0_mask;
  wire [25:0] mem_42_2_R0_addr;
  wire  mem_42_2_R0_clk;
  wire [7:0] mem_42_2_R0_data;
  wire  mem_42_2_R0_en;
  wire [25:0] mem_42_2_W0_addr;
  wire  mem_42_2_W0_clk;
  wire [7:0] mem_42_2_W0_data;
  wire  mem_42_2_W0_en;
  wire  mem_42_2_W0_mask;
  wire [25:0] mem_42_3_R0_addr;
  wire  mem_42_3_R0_clk;
  wire [7:0] mem_42_3_R0_data;
  wire  mem_42_3_R0_en;
  wire [25:0] mem_42_3_W0_addr;
  wire  mem_42_3_W0_clk;
  wire [7:0] mem_42_3_W0_data;
  wire  mem_42_3_W0_en;
  wire  mem_42_3_W0_mask;
  wire [25:0] mem_42_4_R0_addr;
  wire  mem_42_4_R0_clk;
  wire [7:0] mem_42_4_R0_data;
  wire  mem_42_4_R0_en;
  wire [25:0] mem_42_4_W0_addr;
  wire  mem_42_4_W0_clk;
  wire [7:0] mem_42_4_W0_data;
  wire  mem_42_4_W0_en;
  wire  mem_42_4_W0_mask;
  wire [25:0] mem_42_5_R0_addr;
  wire  mem_42_5_R0_clk;
  wire [7:0] mem_42_5_R0_data;
  wire  mem_42_5_R0_en;
  wire [25:0] mem_42_5_W0_addr;
  wire  mem_42_5_W0_clk;
  wire [7:0] mem_42_5_W0_data;
  wire  mem_42_5_W0_en;
  wire  mem_42_5_W0_mask;
  wire [25:0] mem_42_6_R0_addr;
  wire  mem_42_6_R0_clk;
  wire [7:0] mem_42_6_R0_data;
  wire  mem_42_6_R0_en;
  wire [25:0] mem_42_6_W0_addr;
  wire  mem_42_6_W0_clk;
  wire [7:0] mem_42_6_W0_data;
  wire  mem_42_6_W0_en;
  wire  mem_42_6_W0_mask;
  wire [25:0] mem_42_7_R0_addr;
  wire  mem_42_7_R0_clk;
  wire [7:0] mem_42_7_R0_data;
  wire  mem_42_7_R0_en;
  wire [25:0] mem_42_7_W0_addr;
  wire  mem_42_7_W0_clk;
  wire [7:0] mem_42_7_W0_data;
  wire  mem_42_7_W0_en;
  wire  mem_42_7_W0_mask;
  wire [25:0] mem_43_0_R0_addr;
  wire  mem_43_0_R0_clk;
  wire [7:0] mem_43_0_R0_data;
  wire  mem_43_0_R0_en;
  wire [25:0] mem_43_0_W0_addr;
  wire  mem_43_0_W0_clk;
  wire [7:0] mem_43_0_W0_data;
  wire  mem_43_0_W0_en;
  wire  mem_43_0_W0_mask;
  wire [25:0] mem_43_1_R0_addr;
  wire  mem_43_1_R0_clk;
  wire [7:0] mem_43_1_R0_data;
  wire  mem_43_1_R0_en;
  wire [25:0] mem_43_1_W0_addr;
  wire  mem_43_1_W0_clk;
  wire [7:0] mem_43_1_W0_data;
  wire  mem_43_1_W0_en;
  wire  mem_43_1_W0_mask;
  wire [25:0] mem_43_2_R0_addr;
  wire  mem_43_2_R0_clk;
  wire [7:0] mem_43_2_R0_data;
  wire  mem_43_2_R0_en;
  wire [25:0] mem_43_2_W0_addr;
  wire  mem_43_2_W0_clk;
  wire [7:0] mem_43_2_W0_data;
  wire  mem_43_2_W0_en;
  wire  mem_43_2_W0_mask;
  wire [25:0] mem_43_3_R0_addr;
  wire  mem_43_3_R0_clk;
  wire [7:0] mem_43_3_R0_data;
  wire  mem_43_3_R0_en;
  wire [25:0] mem_43_3_W0_addr;
  wire  mem_43_3_W0_clk;
  wire [7:0] mem_43_3_W0_data;
  wire  mem_43_3_W0_en;
  wire  mem_43_3_W0_mask;
  wire [25:0] mem_43_4_R0_addr;
  wire  mem_43_4_R0_clk;
  wire [7:0] mem_43_4_R0_data;
  wire  mem_43_4_R0_en;
  wire [25:0] mem_43_4_W0_addr;
  wire  mem_43_4_W0_clk;
  wire [7:0] mem_43_4_W0_data;
  wire  mem_43_4_W0_en;
  wire  mem_43_4_W0_mask;
  wire [25:0] mem_43_5_R0_addr;
  wire  mem_43_5_R0_clk;
  wire [7:0] mem_43_5_R0_data;
  wire  mem_43_5_R0_en;
  wire [25:0] mem_43_5_W0_addr;
  wire  mem_43_5_W0_clk;
  wire [7:0] mem_43_5_W0_data;
  wire  mem_43_5_W0_en;
  wire  mem_43_5_W0_mask;
  wire [25:0] mem_43_6_R0_addr;
  wire  mem_43_6_R0_clk;
  wire [7:0] mem_43_6_R0_data;
  wire  mem_43_6_R0_en;
  wire [25:0] mem_43_6_W0_addr;
  wire  mem_43_6_W0_clk;
  wire [7:0] mem_43_6_W0_data;
  wire  mem_43_6_W0_en;
  wire  mem_43_6_W0_mask;
  wire [25:0] mem_43_7_R0_addr;
  wire  mem_43_7_R0_clk;
  wire [7:0] mem_43_7_R0_data;
  wire  mem_43_7_R0_en;
  wire [25:0] mem_43_7_W0_addr;
  wire  mem_43_7_W0_clk;
  wire [7:0] mem_43_7_W0_data;
  wire  mem_43_7_W0_en;
  wire  mem_43_7_W0_mask;
  wire [25:0] mem_44_0_R0_addr;
  wire  mem_44_0_R0_clk;
  wire [7:0] mem_44_0_R0_data;
  wire  mem_44_0_R0_en;
  wire [25:0] mem_44_0_W0_addr;
  wire  mem_44_0_W0_clk;
  wire [7:0] mem_44_0_W0_data;
  wire  mem_44_0_W0_en;
  wire  mem_44_0_W0_mask;
  wire [25:0] mem_44_1_R0_addr;
  wire  mem_44_1_R0_clk;
  wire [7:0] mem_44_1_R0_data;
  wire  mem_44_1_R0_en;
  wire [25:0] mem_44_1_W0_addr;
  wire  mem_44_1_W0_clk;
  wire [7:0] mem_44_1_W0_data;
  wire  mem_44_1_W0_en;
  wire  mem_44_1_W0_mask;
  wire [25:0] mem_44_2_R0_addr;
  wire  mem_44_2_R0_clk;
  wire [7:0] mem_44_2_R0_data;
  wire  mem_44_2_R0_en;
  wire [25:0] mem_44_2_W0_addr;
  wire  mem_44_2_W0_clk;
  wire [7:0] mem_44_2_W0_data;
  wire  mem_44_2_W0_en;
  wire  mem_44_2_W0_mask;
  wire [25:0] mem_44_3_R0_addr;
  wire  mem_44_3_R0_clk;
  wire [7:0] mem_44_3_R0_data;
  wire  mem_44_3_R0_en;
  wire [25:0] mem_44_3_W0_addr;
  wire  mem_44_3_W0_clk;
  wire [7:0] mem_44_3_W0_data;
  wire  mem_44_3_W0_en;
  wire  mem_44_3_W0_mask;
  wire [25:0] mem_44_4_R0_addr;
  wire  mem_44_4_R0_clk;
  wire [7:0] mem_44_4_R0_data;
  wire  mem_44_4_R0_en;
  wire [25:0] mem_44_4_W0_addr;
  wire  mem_44_4_W0_clk;
  wire [7:0] mem_44_4_W0_data;
  wire  mem_44_4_W0_en;
  wire  mem_44_4_W0_mask;
  wire [25:0] mem_44_5_R0_addr;
  wire  mem_44_5_R0_clk;
  wire [7:0] mem_44_5_R0_data;
  wire  mem_44_5_R0_en;
  wire [25:0] mem_44_5_W0_addr;
  wire  mem_44_5_W0_clk;
  wire [7:0] mem_44_5_W0_data;
  wire  mem_44_5_W0_en;
  wire  mem_44_5_W0_mask;
  wire [25:0] mem_44_6_R0_addr;
  wire  mem_44_6_R0_clk;
  wire [7:0] mem_44_6_R0_data;
  wire  mem_44_6_R0_en;
  wire [25:0] mem_44_6_W0_addr;
  wire  mem_44_6_W0_clk;
  wire [7:0] mem_44_6_W0_data;
  wire  mem_44_6_W0_en;
  wire  mem_44_6_W0_mask;
  wire [25:0] mem_44_7_R0_addr;
  wire  mem_44_7_R0_clk;
  wire [7:0] mem_44_7_R0_data;
  wire  mem_44_7_R0_en;
  wire [25:0] mem_44_7_W0_addr;
  wire  mem_44_7_W0_clk;
  wire [7:0] mem_44_7_W0_data;
  wire  mem_44_7_W0_en;
  wire  mem_44_7_W0_mask;
  wire [25:0] mem_45_0_R0_addr;
  wire  mem_45_0_R0_clk;
  wire [7:0] mem_45_0_R0_data;
  wire  mem_45_0_R0_en;
  wire [25:0] mem_45_0_W0_addr;
  wire  mem_45_0_W0_clk;
  wire [7:0] mem_45_0_W0_data;
  wire  mem_45_0_W0_en;
  wire  mem_45_0_W0_mask;
  wire [25:0] mem_45_1_R0_addr;
  wire  mem_45_1_R0_clk;
  wire [7:0] mem_45_1_R0_data;
  wire  mem_45_1_R0_en;
  wire [25:0] mem_45_1_W0_addr;
  wire  mem_45_1_W0_clk;
  wire [7:0] mem_45_1_W0_data;
  wire  mem_45_1_W0_en;
  wire  mem_45_1_W0_mask;
  wire [25:0] mem_45_2_R0_addr;
  wire  mem_45_2_R0_clk;
  wire [7:0] mem_45_2_R0_data;
  wire  mem_45_2_R0_en;
  wire [25:0] mem_45_2_W0_addr;
  wire  mem_45_2_W0_clk;
  wire [7:0] mem_45_2_W0_data;
  wire  mem_45_2_W0_en;
  wire  mem_45_2_W0_mask;
  wire [25:0] mem_45_3_R0_addr;
  wire  mem_45_3_R0_clk;
  wire [7:0] mem_45_3_R0_data;
  wire  mem_45_3_R0_en;
  wire [25:0] mem_45_3_W0_addr;
  wire  mem_45_3_W0_clk;
  wire [7:0] mem_45_3_W0_data;
  wire  mem_45_3_W0_en;
  wire  mem_45_3_W0_mask;
  wire [25:0] mem_45_4_R0_addr;
  wire  mem_45_4_R0_clk;
  wire [7:0] mem_45_4_R0_data;
  wire  mem_45_4_R0_en;
  wire [25:0] mem_45_4_W0_addr;
  wire  mem_45_4_W0_clk;
  wire [7:0] mem_45_4_W0_data;
  wire  mem_45_4_W0_en;
  wire  mem_45_4_W0_mask;
  wire [25:0] mem_45_5_R0_addr;
  wire  mem_45_5_R0_clk;
  wire [7:0] mem_45_5_R0_data;
  wire  mem_45_5_R0_en;
  wire [25:0] mem_45_5_W0_addr;
  wire  mem_45_5_W0_clk;
  wire [7:0] mem_45_5_W0_data;
  wire  mem_45_5_W0_en;
  wire  mem_45_5_W0_mask;
  wire [25:0] mem_45_6_R0_addr;
  wire  mem_45_6_R0_clk;
  wire [7:0] mem_45_6_R0_data;
  wire  mem_45_6_R0_en;
  wire [25:0] mem_45_6_W0_addr;
  wire  mem_45_6_W0_clk;
  wire [7:0] mem_45_6_W0_data;
  wire  mem_45_6_W0_en;
  wire  mem_45_6_W0_mask;
  wire [25:0] mem_45_7_R0_addr;
  wire  mem_45_7_R0_clk;
  wire [7:0] mem_45_7_R0_data;
  wire  mem_45_7_R0_en;
  wire [25:0] mem_45_7_W0_addr;
  wire  mem_45_7_W0_clk;
  wire [7:0] mem_45_7_W0_data;
  wire  mem_45_7_W0_en;
  wire  mem_45_7_W0_mask;
  wire [25:0] mem_46_0_R0_addr;
  wire  mem_46_0_R0_clk;
  wire [7:0] mem_46_0_R0_data;
  wire  mem_46_0_R0_en;
  wire [25:0] mem_46_0_W0_addr;
  wire  mem_46_0_W0_clk;
  wire [7:0] mem_46_0_W0_data;
  wire  mem_46_0_W0_en;
  wire  mem_46_0_W0_mask;
  wire [25:0] mem_46_1_R0_addr;
  wire  mem_46_1_R0_clk;
  wire [7:0] mem_46_1_R0_data;
  wire  mem_46_1_R0_en;
  wire [25:0] mem_46_1_W0_addr;
  wire  mem_46_1_W0_clk;
  wire [7:0] mem_46_1_W0_data;
  wire  mem_46_1_W0_en;
  wire  mem_46_1_W0_mask;
  wire [25:0] mem_46_2_R0_addr;
  wire  mem_46_2_R0_clk;
  wire [7:0] mem_46_2_R0_data;
  wire  mem_46_2_R0_en;
  wire [25:0] mem_46_2_W0_addr;
  wire  mem_46_2_W0_clk;
  wire [7:0] mem_46_2_W0_data;
  wire  mem_46_2_W0_en;
  wire  mem_46_2_W0_mask;
  wire [25:0] mem_46_3_R0_addr;
  wire  mem_46_3_R0_clk;
  wire [7:0] mem_46_3_R0_data;
  wire  mem_46_3_R0_en;
  wire [25:0] mem_46_3_W0_addr;
  wire  mem_46_3_W0_clk;
  wire [7:0] mem_46_3_W0_data;
  wire  mem_46_3_W0_en;
  wire  mem_46_3_W0_mask;
  wire [25:0] mem_46_4_R0_addr;
  wire  mem_46_4_R0_clk;
  wire [7:0] mem_46_4_R0_data;
  wire  mem_46_4_R0_en;
  wire [25:0] mem_46_4_W0_addr;
  wire  mem_46_4_W0_clk;
  wire [7:0] mem_46_4_W0_data;
  wire  mem_46_4_W0_en;
  wire  mem_46_4_W0_mask;
  wire [25:0] mem_46_5_R0_addr;
  wire  mem_46_5_R0_clk;
  wire [7:0] mem_46_5_R0_data;
  wire  mem_46_5_R0_en;
  wire [25:0] mem_46_5_W0_addr;
  wire  mem_46_5_W0_clk;
  wire [7:0] mem_46_5_W0_data;
  wire  mem_46_5_W0_en;
  wire  mem_46_5_W0_mask;
  wire [25:0] mem_46_6_R0_addr;
  wire  mem_46_6_R0_clk;
  wire [7:0] mem_46_6_R0_data;
  wire  mem_46_6_R0_en;
  wire [25:0] mem_46_6_W0_addr;
  wire  mem_46_6_W0_clk;
  wire [7:0] mem_46_6_W0_data;
  wire  mem_46_6_W0_en;
  wire  mem_46_6_W0_mask;
  wire [25:0] mem_46_7_R0_addr;
  wire  mem_46_7_R0_clk;
  wire [7:0] mem_46_7_R0_data;
  wire  mem_46_7_R0_en;
  wire [25:0] mem_46_7_W0_addr;
  wire  mem_46_7_W0_clk;
  wire [7:0] mem_46_7_W0_data;
  wire  mem_46_7_W0_en;
  wire  mem_46_7_W0_mask;
  wire [25:0] mem_47_0_R0_addr;
  wire  mem_47_0_R0_clk;
  wire [7:0] mem_47_0_R0_data;
  wire  mem_47_0_R0_en;
  wire [25:0] mem_47_0_W0_addr;
  wire  mem_47_0_W0_clk;
  wire [7:0] mem_47_0_W0_data;
  wire  mem_47_0_W0_en;
  wire  mem_47_0_W0_mask;
  wire [25:0] mem_47_1_R0_addr;
  wire  mem_47_1_R0_clk;
  wire [7:0] mem_47_1_R0_data;
  wire  mem_47_1_R0_en;
  wire [25:0] mem_47_1_W0_addr;
  wire  mem_47_1_W0_clk;
  wire [7:0] mem_47_1_W0_data;
  wire  mem_47_1_W0_en;
  wire  mem_47_1_W0_mask;
  wire [25:0] mem_47_2_R0_addr;
  wire  mem_47_2_R0_clk;
  wire [7:0] mem_47_2_R0_data;
  wire  mem_47_2_R0_en;
  wire [25:0] mem_47_2_W0_addr;
  wire  mem_47_2_W0_clk;
  wire [7:0] mem_47_2_W0_data;
  wire  mem_47_2_W0_en;
  wire  mem_47_2_W0_mask;
  wire [25:0] mem_47_3_R0_addr;
  wire  mem_47_3_R0_clk;
  wire [7:0] mem_47_3_R0_data;
  wire  mem_47_3_R0_en;
  wire [25:0] mem_47_3_W0_addr;
  wire  mem_47_3_W0_clk;
  wire [7:0] mem_47_3_W0_data;
  wire  mem_47_3_W0_en;
  wire  mem_47_3_W0_mask;
  wire [25:0] mem_47_4_R0_addr;
  wire  mem_47_4_R0_clk;
  wire [7:0] mem_47_4_R0_data;
  wire  mem_47_4_R0_en;
  wire [25:0] mem_47_4_W0_addr;
  wire  mem_47_4_W0_clk;
  wire [7:0] mem_47_4_W0_data;
  wire  mem_47_4_W0_en;
  wire  mem_47_4_W0_mask;
  wire [25:0] mem_47_5_R0_addr;
  wire  mem_47_5_R0_clk;
  wire [7:0] mem_47_5_R0_data;
  wire  mem_47_5_R0_en;
  wire [25:0] mem_47_5_W0_addr;
  wire  mem_47_5_W0_clk;
  wire [7:0] mem_47_5_W0_data;
  wire  mem_47_5_W0_en;
  wire  mem_47_5_W0_mask;
  wire [25:0] mem_47_6_R0_addr;
  wire  mem_47_6_R0_clk;
  wire [7:0] mem_47_6_R0_data;
  wire  mem_47_6_R0_en;
  wire [25:0] mem_47_6_W0_addr;
  wire  mem_47_6_W0_clk;
  wire [7:0] mem_47_6_W0_data;
  wire  mem_47_6_W0_en;
  wire  mem_47_6_W0_mask;
  wire [25:0] mem_47_7_R0_addr;
  wire  mem_47_7_R0_clk;
  wire [7:0] mem_47_7_R0_data;
  wire  mem_47_7_R0_en;
  wire [25:0] mem_47_7_W0_addr;
  wire  mem_47_7_W0_clk;
  wire [7:0] mem_47_7_W0_data;
  wire  mem_47_7_W0_en;
  wire  mem_47_7_W0_mask;
  wire [25:0] mem_48_0_R0_addr;
  wire  mem_48_0_R0_clk;
  wire [7:0] mem_48_0_R0_data;
  wire  mem_48_0_R0_en;
  wire [25:0] mem_48_0_W0_addr;
  wire  mem_48_0_W0_clk;
  wire [7:0] mem_48_0_W0_data;
  wire  mem_48_0_W0_en;
  wire  mem_48_0_W0_mask;
  wire [25:0] mem_48_1_R0_addr;
  wire  mem_48_1_R0_clk;
  wire [7:0] mem_48_1_R0_data;
  wire  mem_48_1_R0_en;
  wire [25:0] mem_48_1_W0_addr;
  wire  mem_48_1_W0_clk;
  wire [7:0] mem_48_1_W0_data;
  wire  mem_48_1_W0_en;
  wire  mem_48_1_W0_mask;
  wire [25:0] mem_48_2_R0_addr;
  wire  mem_48_2_R0_clk;
  wire [7:0] mem_48_2_R0_data;
  wire  mem_48_2_R0_en;
  wire [25:0] mem_48_2_W0_addr;
  wire  mem_48_2_W0_clk;
  wire [7:0] mem_48_2_W0_data;
  wire  mem_48_2_W0_en;
  wire  mem_48_2_W0_mask;
  wire [25:0] mem_48_3_R0_addr;
  wire  mem_48_3_R0_clk;
  wire [7:0] mem_48_3_R0_data;
  wire  mem_48_3_R0_en;
  wire [25:0] mem_48_3_W0_addr;
  wire  mem_48_3_W0_clk;
  wire [7:0] mem_48_3_W0_data;
  wire  mem_48_3_W0_en;
  wire  mem_48_3_W0_mask;
  wire [25:0] mem_48_4_R0_addr;
  wire  mem_48_4_R0_clk;
  wire [7:0] mem_48_4_R0_data;
  wire  mem_48_4_R0_en;
  wire [25:0] mem_48_4_W0_addr;
  wire  mem_48_4_W0_clk;
  wire [7:0] mem_48_4_W0_data;
  wire  mem_48_4_W0_en;
  wire  mem_48_4_W0_mask;
  wire [25:0] mem_48_5_R0_addr;
  wire  mem_48_5_R0_clk;
  wire [7:0] mem_48_5_R0_data;
  wire  mem_48_5_R0_en;
  wire [25:0] mem_48_5_W0_addr;
  wire  mem_48_5_W0_clk;
  wire [7:0] mem_48_5_W0_data;
  wire  mem_48_5_W0_en;
  wire  mem_48_5_W0_mask;
  wire [25:0] mem_48_6_R0_addr;
  wire  mem_48_6_R0_clk;
  wire [7:0] mem_48_6_R0_data;
  wire  mem_48_6_R0_en;
  wire [25:0] mem_48_6_W0_addr;
  wire  mem_48_6_W0_clk;
  wire [7:0] mem_48_6_W0_data;
  wire  mem_48_6_W0_en;
  wire  mem_48_6_W0_mask;
  wire [25:0] mem_48_7_R0_addr;
  wire  mem_48_7_R0_clk;
  wire [7:0] mem_48_7_R0_data;
  wire  mem_48_7_R0_en;
  wire [25:0] mem_48_7_W0_addr;
  wire  mem_48_7_W0_clk;
  wire [7:0] mem_48_7_W0_data;
  wire  mem_48_7_W0_en;
  wire  mem_48_7_W0_mask;
  wire [25:0] mem_49_0_R0_addr;
  wire  mem_49_0_R0_clk;
  wire [7:0] mem_49_0_R0_data;
  wire  mem_49_0_R0_en;
  wire [25:0] mem_49_0_W0_addr;
  wire  mem_49_0_W0_clk;
  wire [7:0] mem_49_0_W0_data;
  wire  mem_49_0_W0_en;
  wire  mem_49_0_W0_mask;
  wire [25:0] mem_49_1_R0_addr;
  wire  mem_49_1_R0_clk;
  wire [7:0] mem_49_1_R0_data;
  wire  mem_49_1_R0_en;
  wire [25:0] mem_49_1_W0_addr;
  wire  mem_49_1_W0_clk;
  wire [7:0] mem_49_1_W0_data;
  wire  mem_49_1_W0_en;
  wire  mem_49_1_W0_mask;
  wire [25:0] mem_49_2_R0_addr;
  wire  mem_49_2_R0_clk;
  wire [7:0] mem_49_2_R0_data;
  wire  mem_49_2_R0_en;
  wire [25:0] mem_49_2_W0_addr;
  wire  mem_49_2_W0_clk;
  wire [7:0] mem_49_2_W0_data;
  wire  mem_49_2_W0_en;
  wire  mem_49_2_W0_mask;
  wire [25:0] mem_49_3_R0_addr;
  wire  mem_49_3_R0_clk;
  wire [7:0] mem_49_3_R0_data;
  wire  mem_49_3_R0_en;
  wire [25:0] mem_49_3_W0_addr;
  wire  mem_49_3_W0_clk;
  wire [7:0] mem_49_3_W0_data;
  wire  mem_49_3_W0_en;
  wire  mem_49_3_W0_mask;
  wire [25:0] mem_49_4_R0_addr;
  wire  mem_49_4_R0_clk;
  wire [7:0] mem_49_4_R0_data;
  wire  mem_49_4_R0_en;
  wire [25:0] mem_49_4_W0_addr;
  wire  mem_49_4_W0_clk;
  wire [7:0] mem_49_4_W0_data;
  wire  mem_49_4_W0_en;
  wire  mem_49_4_W0_mask;
  wire [25:0] mem_49_5_R0_addr;
  wire  mem_49_5_R0_clk;
  wire [7:0] mem_49_5_R0_data;
  wire  mem_49_5_R0_en;
  wire [25:0] mem_49_5_W0_addr;
  wire  mem_49_5_W0_clk;
  wire [7:0] mem_49_5_W0_data;
  wire  mem_49_5_W0_en;
  wire  mem_49_5_W0_mask;
  wire [25:0] mem_49_6_R0_addr;
  wire  mem_49_6_R0_clk;
  wire [7:0] mem_49_6_R0_data;
  wire  mem_49_6_R0_en;
  wire [25:0] mem_49_6_W0_addr;
  wire  mem_49_6_W0_clk;
  wire [7:0] mem_49_6_W0_data;
  wire  mem_49_6_W0_en;
  wire  mem_49_6_W0_mask;
  wire [25:0] mem_49_7_R0_addr;
  wire  mem_49_7_R0_clk;
  wire [7:0] mem_49_7_R0_data;
  wire  mem_49_7_R0_en;
  wire [25:0] mem_49_7_W0_addr;
  wire  mem_49_7_W0_clk;
  wire [7:0] mem_49_7_W0_data;
  wire  mem_49_7_W0_en;
  wire  mem_49_7_W0_mask;
  wire [25:0] mem_50_0_R0_addr;
  wire  mem_50_0_R0_clk;
  wire [7:0] mem_50_0_R0_data;
  wire  mem_50_0_R0_en;
  wire [25:0] mem_50_0_W0_addr;
  wire  mem_50_0_W0_clk;
  wire [7:0] mem_50_0_W0_data;
  wire  mem_50_0_W0_en;
  wire  mem_50_0_W0_mask;
  wire [25:0] mem_50_1_R0_addr;
  wire  mem_50_1_R0_clk;
  wire [7:0] mem_50_1_R0_data;
  wire  mem_50_1_R0_en;
  wire [25:0] mem_50_1_W0_addr;
  wire  mem_50_1_W0_clk;
  wire [7:0] mem_50_1_W0_data;
  wire  mem_50_1_W0_en;
  wire  mem_50_1_W0_mask;
  wire [25:0] mem_50_2_R0_addr;
  wire  mem_50_2_R0_clk;
  wire [7:0] mem_50_2_R0_data;
  wire  mem_50_2_R0_en;
  wire [25:0] mem_50_2_W0_addr;
  wire  mem_50_2_W0_clk;
  wire [7:0] mem_50_2_W0_data;
  wire  mem_50_2_W0_en;
  wire  mem_50_2_W0_mask;
  wire [25:0] mem_50_3_R0_addr;
  wire  mem_50_3_R0_clk;
  wire [7:0] mem_50_3_R0_data;
  wire  mem_50_3_R0_en;
  wire [25:0] mem_50_3_W0_addr;
  wire  mem_50_3_W0_clk;
  wire [7:0] mem_50_3_W0_data;
  wire  mem_50_3_W0_en;
  wire  mem_50_3_W0_mask;
  wire [25:0] mem_50_4_R0_addr;
  wire  mem_50_4_R0_clk;
  wire [7:0] mem_50_4_R0_data;
  wire  mem_50_4_R0_en;
  wire [25:0] mem_50_4_W0_addr;
  wire  mem_50_4_W0_clk;
  wire [7:0] mem_50_4_W0_data;
  wire  mem_50_4_W0_en;
  wire  mem_50_4_W0_mask;
  wire [25:0] mem_50_5_R0_addr;
  wire  mem_50_5_R0_clk;
  wire [7:0] mem_50_5_R0_data;
  wire  mem_50_5_R0_en;
  wire [25:0] mem_50_5_W0_addr;
  wire  mem_50_5_W0_clk;
  wire [7:0] mem_50_5_W0_data;
  wire  mem_50_5_W0_en;
  wire  mem_50_5_W0_mask;
  wire [25:0] mem_50_6_R0_addr;
  wire  mem_50_6_R0_clk;
  wire [7:0] mem_50_6_R0_data;
  wire  mem_50_6_R0_en;
  wire [25:0] mem_50_6_W0_addr;
  wire  mem_50_6_W0_clk;
  wire [7:0] mem_50_6_W0_data;
  wire  mem_50_6_W0_en;
  wire  mem_50_6_W0_mask;
  wire [25:0] mem_50_7_R0_addr;
  wire  mem_50_7_R0_clk;
  wire [7:0] mem_50_7_R0_data;
  wire  mem_50_7_R0_en;
  wire [25:0] mem_50_7_W0_addr;
  wire  mem_50_7_W0_clk;
  wire [7:0] mem_50_7_W0_data;
  wire  mem_50_7_W0_en;
  wire  mem_50_7_W0_mask;
  wire [25:0] mem_51_0_R0_addr;
  wire  mem_51_0_R0_clk;
  wire [7:0] mem_51_0_R0_data;
  wire  mem_51_0_R0_en;
  wire [25:0] mem_51_0_W0_addr;
  wire  mem_51_0_W0_clk;
  wire [7:0] mem_51_0_W0_data;
  wire  mem_51_0_W0_en;
  wire  mem_51_0_W0_mask;
  wire [25:0] mem_51_1_R0_addr;
  wire  mem_51_1_R0_clk;
  wire [7:0] mem_51_1_R0_data;
  wire  mem_51_1_R0_en;
  wire [25:0] mem_51_1_W0_addr;
  wire  mem_51_1_W0_clk;
  wire [7:0] mem_51_1_W0_data;
  wire  mem_51_1_W0_en;
  wire  mem_51_1_W0_mask;
  wire [25:0] mem_51_2_R0_addr;
  wire  mem_51_2_R0_clk;
  wire [7:0] mem_51_2_R0_data;
  wire  mem_51_2_R0_en;
  wire [25:0] mem_51_2_W0_addr;
  wire  mem_51_2_W0_clk;
  wire [7:0] mem_51_2_W0_data;
  wire  mem_51_2_W0_en;
  wire  mem_51_2_W0_mask;
  wire [25:0] mem_51_3_R0_addr;
  wire  mem_51_3_R0_clk;
  wire [7:0] mem_51_3_R0_data;
  wire  mem_51_3_R0_en;
  wire [25:0] mem_51_3_W0_addr;
  wire  mem_51_3_W0_clk;
  wire [7:0] mem_51_3_W0_data;
  wire  mem_51_3_W0_en;
  wire  mem_51_3_W0_mask;
  wire [25:0] mem_51_4_R0_addr;
  wire  mem_51_4_R0_clk;
  wire [7:0] mem_51_4_R0_data;
  wire  mem_51_4_R0_en;
  wire [25:0] mem_51_4_W0_addr;
  wire  mem_51_4_W0_clk;
  wire [7:0] mem_51_4_W0_data;
  wire  mem_51_4_W0_en;
  wire  mem_51_4_W0_mask;
  wire [25:0] mem_51_5_R0_addr;
  wire  mem_51_5_R0_clk;
  wire [7:0] mem_51_5_R0_data;
  wire  mem_51_5_R0_en;
  wire [25:0] mem_51_5_W0_addr;
  wire  mem_51_5_W0_clk;
  wire [7:0] mem_51_5_W0_data;
  wire  mem_51_5_W0_en;
  wire  mem_51_5_W0_mask;
  wire [25:0] mem_51_6_R0_addr;
  wire  mem_51_6_R0_clk;
  wire [7:0] mem_51_6_R0_data;
  wire  mem_51_6_R0_en;
  wire [25:0] mem_51_6_W0_addr;
  wire  mem_51_6_W0_clk;
  wire [7:0] mem_51_6_W0_data;
  wire  mem_51_6_W0_en;
  wire  mem_51_6_W0_mask;
  wire [25:0] mem_51_7_R0_addr;
  wire  mem_51_7_R0_clk;
  wire [7:0] mem_51_7_R0_data;
  wire  mem_51_7_R0_en;
  wire [25:0] mem_51_7_W0_addr;
  wire  mem_51_7_W0_clk;
  wire [7:0] mem_51_7_W0_data;
  wire  mem_51_7_W0_en;
  wire  mem_51_7_W0_mask;
  wire [25:0] mem_52_0_R0_addr;
  wire  mem_52_0_R0_clk;
  wire [7:0] mem_52_0_R0_data;
  wire  mem_52_0_R0_en;
  wire [25:0] mem_52_0_W0_addr;
  wire  mem_52_0_W0_clk;
  wire [7:0] mem_52_0_W0_data;
  wire  mem_52_0_W0_en;
  wire  mem_52_0_W0_mask;
  wire [25:0] mem_52_1_R0_addr;
  wire  mem_52_1_R0_clk;
  wire [7:0] mem_52_1_R0_data;
  wire  mem_52_1_R0_en;
  wire [25:0] mem_52_1_W0_addr;
  wire  mem_52_1_W0_clk;
  wire [7:0] mem_52_1_W0_data;
  wire  mem_52_1_W0_en;
  wire  mem_52_1_W0_mask;
  wire [25:0] mem_52_2_R0_addr;
  wire  mem_52_2_R0_clk;
  wire [7:0] mem_52_2_R0_data;
  wire  mem_52_2_R0_en;
  wire [25:0] mem_52_2_W0_addr;
  wire  mem_52_2_W0_clk;
  wire [7:0] mem_52_2_W0_data;
  wire  mem_52_2_W0_en;
  wire  mem_52_2_W0_mask;
  wire [25:0] mem_52_3_R0_addr;
  wire  mem_52_3_R0_clk;
  wire [7:0] mem_52_3_R0_data;
  wire  mem_52_3_R0_en;
  wire [25:0] mem_52_3_W0_addr;
  wire  mem_52_3_W0_clk;
  wire [7:0] mem_52_3_W0_data;
  wire  mem_52_3_W0_en;
  wire  mem_52_3_W0_mask;
  wire [25:0] mem_52_4_R0_addr;
  wire  mem_52_4_R0_clk;
  wire [7:0] mem_52_4_R0_data;
  wire  mem_52_4_R0_en;
  wire [25:0] mem_52_4_W0_addr;
  wire  mem_52_4_W0_clk;
  wire [7:0] mem_52_4_W0_data;
  wire  mem_52_4_W0_en;
  wire  mem_52_4_W0_mask;
  wire [25:0] mem_52_5_R0_addr;
  wire  mem_52_5_R0_clk;
  wire [7:0] mem_52_5_R0_data;
  wire  mem_52_5_R0_en;
  wire [25:0] mem_52_5_W0_addr;
  wire  mem_52_5_W0_clk;
  wire [7:0] mem_52_5_W0_data;
  wire  mem_52_5_W0_en;
  wire  mem_52_5_W0_mask;
  wire [25:0] mem_52_6_R0_addr;
  wire  mem_52_6_R0_clk;
  wire [7:0] mem_52_6_R0_data;
  wire  mem_52_6_R0_en;
  wire [25:0] mem_52_6_W0_addr;
  wire  mem_52_6_W0_clk;
  wire [7:0] mem_52_6_W0_data;
  wire  mem_52_6_W0_en;
  wire  mem_52_6_W0_mask;
  wire [25:0] mem_52_7_R0_addr;
  wire  mem_52_7_R0_clk;
  wire [7:0] mem_52_7_R0_data;
  wire  mem_52_7_R0_en;
  wire [25:0] mem_52_7_W0_addr;
  wire  mem_52_7_W0_clk;
  wire [7:0] mem_52_7_W0_data;
  wire  mem_52_7_W0_en;
  wire  mem_52_7_W0_mask;
  wire [25:0] mem_53_0_R0_addr;
  wire  mem_53_0_R0_clk;
  wire [7:0] mem_53_0_R0_data;
  wire  mem_53_0_R0_en;
  wire [25:0] mem_53_0_W0_addr;
  wire  mem_53_0_W0_clk;
  wire [7:0] mem_53_0_W0_data;
  wire  mem_53_0_W0_en;
  wire  mem_53_0_W0_mask;
  wire [25:0] mem_53_1_R0_addr;
  wire  mem_53_1_R0_clk;
  wire [7:0] mem_53_1_R0_data;
  wire  mem_53_1_R0_en;
  wire [25:0] mem_53_1_W0_addr;
  wire  mem_53_1_W0_clk;
  wire [7:0] mem_53_1_W0_data;
  wire  mem_53_1_W0_en;
  wire  mem_53_1_W0_mask;
  wire [25:0] mem_53_2_R0_addr;
  wire  mem_53_2_R0_clk;
  wire [7:0] mem_53_2_R0_data;
  wire  mem_53_2_R0_en;
  wire [25:0] mem_53_2_W0_addr;
  wire  mem_53_2_W0_clk;
  wire [7:0] mem_53_2_W0_data;
  wire  mem_53_2_W0_en;
  wire  mem_53_2_W0_mask;
  wire [25:0] mem_53_3_R0_addr;
  wire  mem_53_3_R0_clk;
  wire [7:0] mem_53_3_R0_data;
  wire  mem_53_3_R0_en;
  wire [25:0] mem_53_3_W0_addr;
  wire  mem_53_3_W0_clk;
  wire [7:0] mem_53_3_W0_data;
  wire  mem_53_3_W0_en;
  wire  mem_53_3_W0_mask;
  wire [25:0] mem_53_4_R0_addr;
  wire  mem_53_4_R0_clk;
  wire [7:0] mem_53_4_R0_data;
  wire  mem_53_4_R0_en;
  wire [25:0] mem_53_4_W0_addr;
  wire  mem_53_4_W0_clk;
  wire [7:0] mem_53_4_W0_data;
  wire  mem_53_4_W0_en;
  wire  mem_53_4_W0_mask;
  wire [25:0] mem_53_5_R0_addr;
  wire  mem_53_5_R0_clk;
  wire [7:0] mem_53_5_R0_data;
  wire  mem_53_5_R0_en;
  wire [25:0] mem_53_5_W0_addr;
  wire  mem_53_5_W0_clk;
  wire [7:0] mem_53_5_W0_data;
  wire  mem_53_5_W0_en;
  wire  mem_53_5_W0_mask;
  wire [25:0] mem_53_6_R0_addr;
  wire  mem_53_6_R0_clk;
  wire [7:0] mem_53_6_R0_data;
  wire  mem_53_6_R0_en;
  wire [25:0] mem_53_6_W0_addr;
  wire  mem_53_6_W0_clk;
  wire [7:0] mem_53_6_W0_data;
  wire  mem_53_6_W0_en;
  wire  mem_53_6_W0_mask;
  wire [25:0] mem_53_7_R0_addr;
  wire  mem_53_7_R0_clk;
  wire [7:0] mem_53_7_R0_data;
  wire  mem_53_7_R0_en;
  wire [25:0] mem_53_7_W0_addr;
  wire  mem_53_7_W0_clk;
  wire [7:0] mem_53_7_W0_data;
  wire  mem_53_7_W0_en;
  wire  mem_53_7_W0_mask;
  wire [25:0] mem_54_0_R0_addr;
  wire  mem_54_0_R0_clk;
  wire [7:0] mem_54_0_R0_data;
  wire  mem_54_0_R0_en;
  wire [25:0] mem_54_0_W0_addr;
  wire  mem_54_0_W0_clk;
  wire [7:0] mem_54_0_W0_data;
  wire  mem_54_0_W0_en;
  wire  mem_54_0_W0_mask;
  wire [25:0] mem_54_1_R0_addr;
  wire  mem_54_1_R0_clk;
  wire [7:0] mem_54_1_R0_data;
  wire  mem_54_1_R0_en;
  wire [25:0] mem_54_1_W0_addr;
  wire  mem_54_1_W0_clk;
  wire [7:0] mem_54_1_W0_data;
  wire  mem_54_1_W0_en;
  wire  mem_54_1_W0_mask;
  wire [25:0] mem_54_2_R0_addr;
  wire  mem_54_2_R0_clk;
  wire [7:0] mem_54_2_R0_data;
  wire  mem_54_2_R0_en;
  wire [25:0] mem_54_2_W0_addr;
  wire  mem_54_2_W0_clk;
  wire [7:0] mem_54_2_W0_data;
  wire  mem_54_2_W0_en;
  wire  mem_54_2_W0_mask;
  wire [25:0] mem_54_3_R0_addr;
  wire  mem_54_3_R0_clk;
  wire [7:0] mem_54_3_R0_data;
  wire  mem_54_3_R0_en;
  wire [25:0] mem_54_3_W0_addr;
  wire  mem_54_3_W0_clk;
  wire [7:0] mem_54_3_W0_data;
  wire  mem_54_3_W0_en;
  wire  mem_54_3_W0_mask;
  wire [25:0] mem_54_4_R0_addr;
  wire  mem_54_4_R0_clk;
  wire [7:0] mem_54_4_R0_data;
  wire  mem_54_4_R0_en;
  wire [25:0] mem_54_4_W0_addr;
  wire  mem_54_4_W0_clk;
  wire [7:0] mem_54_4_W0_data;
  wire  mem_54_4_W0_en;
  wire  mem_54_4_W0_mask;
  wire [25:0] mem_54_5_R0_addr;
  wire  mem_54_5_R0_clk;
  wire [7:0] mem_54_5_R0_data;
  wire  mem_54_5_R0_en;
  wire [25:0] mem_54_5_W0_addr;
  wire  mem_54_5_W0_clk;
  wire [7:0] mem_54_5_W0_data;
  wire  mem_54_5_W0_en;
  wire  mem_54_5_W0_mask;
  wire [25:0] mem_54_6_R0_addr;
  wire  mem_54_6_R0_clk;
  wire [7:0] mem_54_6_R0_data;
  wire  mem_54_6_R0_en;
  wire [25:0] mem_54_6_W0_addr;
  wire  mem_54_6_W0_clk;
  wire [7:0] mem_54_6_W0_data;
  wire  mem_54_6_W0_en;
  wire  mem_54_6_W0_mask;
  wire [25:0] mem_54_7_R0_addr;
  wire  mem_54_7_R0_clk;
  wire [7:0] mem_54_7_R0_data;
  wire  mem_54_7_R0_en;
  wire [25:0] mem_54_7_W0_addr;
  wire  mem_54_7_W0_clk;
  wire [7:0] mem_54_7_W0_data;
  wire  mem_54_7_W0_en;
  wire  mem_54_7_W0_mask;
  wire [25:0] mem_55_0_R0_addr;
  wire  mem_55_0_R0_clk;
  wire [7:0] mem_55_0_R0_data;
  wire  mem_55_0_R0_en;
  wire [25:0] mem_55_0_W0_addr;
  wire  mem_55_0_W0_clk;
  wire [7:0] mem_55_0_W0_data;
  wire  mem_55_0_W0_en;
  wire  mem_55_0_W0_mask;
  wire [25:0] mem_55_1_R0_addr;
  wire  mem_55_1_R0_clk;
  wire [7:0] mem_55_1_R0_data;
  wire  mem_55_1_R0_en;
  wire [25:0] mem_55_1_W0_addr;
  wire  mem_55_1_W0_clk;
  wire [7:0] mem_55_1_W0_data;
  wire  mem_55_1_W0_en;
  wire  mem_55_1_W0_mask;
  wire [25:0] mem_55_2_R0_addr;
  wire  mem_55_2_R0_clk;
  wire [7:0] mem_55_2_R0_data;
  wire  mem_55_2_R0_en;
  wire [25:0] mem_55_2_W0_addr;
  wire  mem_55_2_W0_clk;
  wire [7:0] mem_55_2_W0_data;
  wire  mem_55_2_W0_en;
  wire  mem_55_2_W0_mask;
  wire [25:0] mem_55_3_R0_addr;
  wire  mem_55_3_R0_clk;
  wire [7:0] mem_55_3_R0_data;
  wire  mem_55_3_R0_en;
  wire [25:0] mem_55_3_W0_addr;
  wire  mem_55_3_W0_clk;
  wire [7:0] mem_55_3_W0_data;
  wire  mem_55_3_W0_en;
  wire  mem_55_3_W0_mask;
  wire [25:0] mem_55_4_R0_addr;
  wire  mem_55_4_R0_clk;
  wire [7:0] mem_55_4_R0_data;
  wire  mem_55_4_R0_en;
  wire [25:0] mem_55_4_W0_addr;
  wire  mem_55_4_W0_clk;
  wire [7:0] mem_55_4_W0_data;
  wire  mem_55_4_W0_en;
  wire  mem_55_4_W0_mask;
  wire [25:0] mem_55_5_R0_addr;
  wire  mem_55_5_R0_clk;
  wire [7:0] mem_55_5_R0_data;
  wire  mem_55_5_R0_en;
  wire [25:0] mem_55_5_W0_addr;
  wire  mem_55_5_W0_clk;
  wire [7:0] mem_55_5_W0_data;
  wire  mem_55_5_W0_en;
  wire  mem_55_5_W0_mask;
  wire [25:0] mem_55_6_R0_addr;
  wire  mem_55_6_R0_clk;
  wire [7:0] mem_55_6_R0_data;
  wire  mem_55_6_R0_en;
  wire [25:0] mem_55_6_W0_addr;
  wire  mem_55_6_W0_clk;
  wire [7:0] mem_55_6_W0_data;
  wire  mem_55_6_W0_en;
  wire  mem_55_6_W0_mask;
  wire [25:0] mem_55_7_R0_addr;
  wire  mem_55_7_R0_clk;
  wire [7:0] mem_55_7_R0_data;
  wire  mem_55_7_R0_en;
  wire [25:0] mem_55_7_W0_addr;
  wire  mem_55_7_W0_clk;
  wire [7:0] mem_55_7_W0_data;
  wire  mem_55_7_W0_en;
  wire  mem_55_7_W0_mask;
  wire [25:0] mem_56_0_R0_addr;
  wire  mem_56_0_R0_clk;
  wire [7:0] mem_56_0_R0_data;
  wire  mem_56_0_R0_en;
  wire [25:0] mem_56_0_W0_addr;
  wire  mem_56_0_W0_clk;
  wire [7:0] mem_56_0_W0_data;
  wire  mem_56_0_W0_en;
  wire  mem_56_0_W0_mask;
  wire [25:0] mem_56_1_R0_addr;
  wire  mem_56_1_R0_clk;
  wire [7:0] mem_56_1_R0_data;
  wire  mem_56_1_R0_en;
  wire [25:0] mem_56_1_W0_addr;
  wire  mem_56_1_W0_clk;
  wire [7:0] mem_56_1_W0_data;
  wire  mem_56_1_W0_en;
  wire  mem_56_1_W0_mask;
  wire [25:0] mem_56_2_R0_addr;
  wire  mem_56_2_R0_clk;
  wire [7:0] mem_56_2_R0_data;
  wire  mem_56_2_R0_en;
  wire [25:0] mem_56_2_W0_addr;
  wire  mem_56_2_W0_clk;
  wire [7:0] mem_56_2_W0_data;
  wire  mem_56_2_W0_en;
  wire  mem_56_2_W0_mask;
  wire [25:0] mem_56_3_R0_addr;
  wire  mem_56_3_R0_clk;
  wire [7:0] mem_56_3_R0_data;
  wire  mem_56_3_R0_en;
  wire [25:0] mem_56_3_W0_addr;
  wire  mem_56_3_W0_clk;
  wire [7:0] mem_56_3_W0_data;
  wire  mem_56_3_W0_en;
  wire  mem_56_3_W0_mask;
  wire [25:0] mem_56_4_R0_addr;
  wire  mem_56_4_R0_clk;
  wire [7:0] mem_56_4_R0_data;
  wire  mem_56_4_R0_en;
  wire [25:0] mem_56_4_W0_addr;
  wire  mem_56_4_W0_clk;
  wire [7:0] mem_56_4_W0_data;
  wire  mem_56_4_W0_en;
  wire  mem_56_4_W0_mask;
  wire [25:0] mem_56_5_R0_addr;
  wire  mem_56_5_R0_clk;
  wire [7:0] mem_56_5_R0_data;
  wire  mem_56_5_R0_en;
  wire [25:0] mem_56_5_W0_addr;
  wire  mem_56_5_W0_clk;
  wire [7:0] mem_56_5_W0_data;
  wire  mem_56_5_W0_en;
  wire  mem_56_5_W0_mask;
  wire [25:0] mem_56_6_R0_addr;
  wire  mem_56_6_R0_clk;
  wire [7:0] mem_56_6_R0_data;
  wire  mem_56_6_R0_en;
  wire [25:0] mem_56_6_W0_addr;
  wire  mem_56_6_W0_clk;
  wire [7:0] mem_56_6_W0_data;
  wire  mem_56_6_W0_en;
  wire  mem_56_6_W0_mask;
  wire [25:0] mem_56_7_R0_addr;
  wire  mem_56_7_R0_clk;
  wire [7:0] mem_56_7_R0_data;
  wire  mem_56_7_R0_en;
  wire [25:0] mem_56_7_W0_addr;
  wire  mem_56_7_W0_clk;
  wire [7:0] mem_56_7_W0_data;
  wire  mem_56_7_W0_en;
  wire  mem_56_7_W0_mask;
  wire [25:0] mem_57_0_R0_addr;
  wire  mem_57_0_R0_clk;
  wire [7:0] mem_57_0_R0_data;
  wire  mem_57_0_R0_en;
  wire [25:0] mem_57_0_W0_addr;
  wire  mem_57_0_W0_clk;
  wire [7:0] mem_57_0_W0_data;
  wire  mem_57_0_W0_en;
  wire  mem_57_0_W0_mask;
  wire [25:0] mem_57_1_R0_addr;
  wire  mem_57_1_R0_clk;
  wire [7:0] mem_57_1_R0_data;
  wire  mem_57_1_R0_en;
  wire [25:0] mem_57_1_W0_addr;
  wire  mem_57_1_W0_clk;
  wire [7:0] mem_57_1_W0_data;
  wire  mem_57_1_W0_en;
  wire  mem_57_1_W0_mask;
  wire [25:0] mem_57_2_R0_addr;
  wire  mem_57_2_R0_clk;
  wire [7:0] mem_57_2_R0_data;
  wire  mem_57_2_R0_en;
  wire [25:0] mem_57_2_W0_addr;
  wire  mem_57_2_W0_clk;
  wire [7:0] mem_57_2_W0_data;
  wire  mem_57_2_W0_en;
  wire  mem_57_2_W0_mask;
  wire [25:0] mem_57_3_R0_addr;
  wire  mem_57_3_R0_clk;
  wire [7:0] mem_57_3_R0_data;
  wire  mem_57_3_R0_en;
  wire [25:0] mem_57_3_W0_addr;
  wire  mem_57_3_W0_clk;
  wire [7:0] mem_57_3_W0_data;
  wire  mem_57_3_W0_en;
  wire  mem_57_3_W0_mask;
  wire [25:0] mem_57_4_R0_addr;
  wire  mem_57_4_R0_clk;
  wire [7:0] mem_57_4_R0_data;
  wire  mem_57_4_R0_en;
  wire [25:0] mem_57_4_W0_addr;
  wire  mem_57_4_W0_clk;
  wire [7:0] mem_57_4_W0_data;
  wire  mem_57_4_W0_en;
  wire  mem_57_4_W0_mask;
  wire [25:0] mem_57_5_R0_addr;
  wire  mem_57_5_R0_clk;
  wire [7:0] mem_57_5_R0_data;
  wire  mem_57_5_R0_en;
  wire [25:0] mem_57_5_W0_addr;
  wire  mem_57_5_W0_clk;
  wire [7:0] mem_57_5_W0_data;
  wire  mem_57_5_W0_en;
  wire  mem_57_5_W0_mask;
  wire [25:0] mem_57_6_R0_addr;
  wire  mem_57_6_R0_clk;
  wire [7:0] mem_57_6_R0_data;
  wire  mem_57_6_R0_en;
  wire [25:0] mem_57_6_W0_addr;
  wire  mem_57_6_W0_clk;
  wire [7:0] mem_57_6_W0_data;
  wire  mem_57_6_W0_en;
  wire  mem_57_6_W0_mask;
  wire [25:0] mem_57_7_R0_addr;
  wire  mem_57_7_R0_clk;
  wire [7:0] mem_57_7_R0_data;
  wire  mem_57_7_R0_en;
  wire [25:0] mem_57_7_W0_addr;
  wire  mem_57_7_W0_clk;
  wire [7:0] mem_57_7_W0_data;
  wire  mem_57_7_W0_en;
  wire  mem_57_7_W0_mask;
  wire [25:0] mem_58_0_R0_addr;
  wire  mem_58_0_R0_clk;
  wire [7:0] mem_58_0_R0_data;
  wire  mem_58_0_R0_en;
  wire [25:0] mem_58_0_W0_addr;
  wire  mem_58_0_W0_clk;
  wire [7:0] mem_58_0_W0_data;
  wire  mem_58_0_W0_en;
  wire  mem_58_0_W0_mask;
  wire [25:0] mem_58_1_R0_addr;
  wire  mem_58_1_R0_clk;
  wire [7:0] mem_58_1_R0_data;
  wire  mem_58_1_R0_en;
  wire [25:0] mem_58_1_W0_addr;
  wire  mem_58_1_W0_clk;
  wire [7:0] mem_58_1_W0_data;
  wire  mem_58_1_W0_en;
  wire  mem_58_1_W0_mask;
  wire [25:0] mem_58_2_R0_addr;
  wire  mem_58_2_R0_clk;
  wire [7:0] mem_58_2_R0_data;
  wire  mem_58_2_R0_en;
  wire [25:0] mem_58_2_W0_addr;
  wire  mem_58_2_W0_clk;
  wire [7:0] mem_58_2_W0_data;
  wire  mem_58_2_W0_en;
  wire  mem_58_2_W0_mask;
  wire [25:0] mem_58_3_R0_addr;
  wire  mem_58_3_R0_clk;
  wire [7:0] mem_58_3_R0_data;
  wire  mem_58_3_R0_en;
  wire [25:0] mem_58_3_W0_addr;
  wire  mem_58_3_W0_clk;
  wire [7:0] mem_58_3_W0_data;
  wire  mem_58_3_W0_en;
  wire  mem_58_3_W0_mask;
  wire [25:0] mem_58_4_R0_addr;
  wire  mem_58_4_R0_clk;
  wire [7:0] mem_58_4_R0_data;
  wire  mem_58_4_R0_en;
  wire [25:0] mem_58_4_W0_addr;
  wire  mem_58_4_W0_clk;
  wire [7:0] mem_58_4_W0_data;
  wire  mem_58_4_W0_en;
  wire  mem_58_4_W0_mask;
  wire [25:0] mem_58_5_R0_addr;
  wire  mem_58_5_R0_clk;
  wire [7:0] mem_58_5_R0_data;
  wire  mem_58_5_R0_en;
  wire [25:0] mem_58_5_W0_addr;
  wire  mem_58_5_W0_clk;
  wire [7:0] mem_58_5_W0_data;
  wire  mem_58_5_W0_en;
  wire  mem_58_5_W0_mask;
  wire [25:0] mem_58_6_R0_addr;
  wire  mem_58_6_R0_clk;
  wire [7:0] mem_58_6_R0_data;
  wire  mem_58_6_R0_en;
  wire [25:0] mem_58_6_W0_addr;
  wire  mem_58_6_W0_clk;
  wire [7:0] mem_58_6_W0_data;
  wire  mem_58_6_W0_en;
  wire  mem_58_6_W0_mask;
  wire [25:0] mem_58_7_R0_addr;
  wire  mem_58_7_R0_clk;
  wire [7:0] mem_58_7_R0_data;
  wire  mem_58_7_R0_en;
  wire [25:0] mem_58_7_W0_addr;
  wire  mem_58_7_W0_clk;
  wire [7:0] mem_58_7_W0_data;
  wire  mem_58_7_W0_en;
  wire  mem_58_7_W0_mask;
  wire [25:0] mem_59_0_R0_addr;
  wire  mem_59_0_R0_clk;
  wire [7:0] mem_59_0_R0_data;
  wire  mem_59_0_R0_en;
  wire [25:0] mem_59_0_W0_addr;
  wire  mem_59_0_W0_clk;
  wire [7:0] mem_59_0_W0_data;
  wire  mem_59_0_W0_en;
  wire  mem_59_0_W0_mask;
  wire [25:0] mem_59_1_R0_addr;
  wire  mem_59_1_R0_clk;
  wire [7:0] mem_59_1_R0_data;
  wire  mem_59_1_R0_en;
  wire [25:0] mem_59_1_W0_addr;
  wire  mem_59_1_W0_clk;
  wire [7:0] mem_59_1_W0_data;
  wire  mem_59_1_W0_en;
  wire  mem_59_1_W0_mask;
  wire [25:0] mem_59_2_R0_addr;
  wire  mem_59_2_R0_clk;
  wire [7:0] mem_59_2_R0_data;
  wire  mem_59_2_R0_en;
  wire [25:0] mem_59_2_W0_addr;
  wire  mem_59_2_W0_clk;
  wire [7:0] mem_59_2_W0_data;
  wire  mem_59_2_W0_en;
  wire  mem_59_2_W0_mask;
  wire [25:0] mem_59_3_R0_addr;
  wire  mem_59_3_R0_clk;
  wire [7:0] mem_59_3_R0_data;
  wire  mem_59_3_R0_en;
  wire [25:0] mem_59_3_W0_addr;
  wire  mem_59_3_W0_clk;
  wire [7:0] mem_59_3_W0_data;
  wire  mem_59_3_W0_en;
  wire  mem_59_3_W0_mask;
  wire [25:0] mem_59_4_R0_addr;
  wire  mem_59_4_R0_clk;
  wire [7:0] mem_59_4_R0_data;
  wire  mem_59_4_R0_en;
  wire [25:0] mem_59_4_W0_addr;
  wire  mem_59_4_W0_clk;
  wire [7:0] mem_59_4_W0_data;
  wire  mem_59_4_W0_en;
  wire  mem_59_4_W0_mask;
  wire [25:0] mem_59_5_R0_addr;
  wire  mem_59_5_R0_clk;
  wire [7:0] mem_59_5_R0_data;
  wire  mem_59_5_R0_en;
  wire [25:0] mem_59_5_W0_addr;
  wire  mem_59_5_W0_clk;
  wire [7:0] mem_59_5_W0_data;
  wire  mem_59_5_W0_en;
  wire  mem_59_5_W0_mask;
  wire [25:0] mem_59_6_R0_addr;
  wire  mem_59_6_R0_clk;
  wire [7:0] mem_59_6_R0_data;
  wire  mem_59_6_R0_en;
  wire [25:0] mem_59_6_W0_addr;
  wire  mem_59_6_W0_clk;
  wire [7:0] mem_59_6_W0_data;
  wire  mem_59_6_W0_en;
  wire  mem_59_6_W0_mask;
  wire [25:0] mem_59_7_R0_addr;
  wire  mem_59_7_R0_clk;
  wire [7:0] mem_59_7_R0_data;
  wire  mem_59_7_R0_en;
  wire [25:0] mem_59_7_W0_addr;
  wire  mem_59_7_W0_clk;
  wire [7:0] mem_59_7_W0_data;
  wire  mem_59_7_W0_en;
  wire  mem_59_7_W0_mask;
  wire [25:0] mem_60_0_R0_addr;
  wire  mem_60_0_R0_clk;
  wire [7:0] mem_60_0_R0_data;
  wire  mem_60_0_R0_en;
  wire [25:0] mem_60_0_W0_addr;
  wire  mem_60_0_W0_clk;
  wire [7:0] mem_60_0_W0_data;
  wire  mem_60_0_W0_en;
  wire  mem_60_0_W0_mask;
  wire [25:0] mem_60_1_R0_addr;
  wire  mem_60_1_R0_clk;
  wire [7:0] mem_60_1_R0_data;
  wire  mem_60_1_R0_en;
  wire [25:0] mem_60_1_W0_addr;
  wire  mem_60_1_W0_clk;
  wire [7:0] mem_60_1_W0_data;
  wire  mem_60_1_W0_en;
  wire  mem_60_1_W0_mask;
  wire [25:0] mem_60_2_R0_addr;
  wire  mem_60_2_R0_clk;
  wire [7:0] mem_60_2_R0_data;
  wire  mem_60_2_R0_en;
  wire [25:0] mem_60_2_W0_addr;
  wire  mem_60_2_W0_clk;
  wire [7:0] mem_60_2_W0_data;
  wire  mem_60_2_W0_en;
  wire  mem_60_2_W0_mask;
  wire [25:0] mem_60_3_R0_addr;
  wire  mem_60_3_R0_clk;
  wire [7:0] mem_60_3_R0_data;
  wire  mem_60_3_R0_en;
  wire [25:0] mem_60_3_W0_addr;
  wire  mem_60_3_W0_clk;
  wire [7:0] mem_60_3_W0_data;
  wire  mem_60_3_W0_en;
  wire  mem_60_3_W0_mask;
  wire [25:0] mem_60_4_R0_addr;
  wire  mem_60_4_R0_clk;
  wire [7:0] mem_60_4_R0_data;
  wire  mem_60_4_R0_en;
  wire [25:0] mem_60_4_W0_addr;
  wire  mem_60_4_W0_clk;
  wire [7:0] mem_60_4_W0_data;
  wire  mem_60_4_W0_en;
  wire  mem_60_4_W0_mask;
  wire [25:0] mem_60_5_R0_addr;
  wire  mem_60_5_R0_clk;
  wire [7:0] mem_60_5_R0_data;
  wire  mem_60_5_R0_en;
  wire [25:0] mem_60_5_W0_addr;
  wire  mem_60_5_W0_clk;
  wire [7:0] mem_60_5_W0_data;
  wire  mem_60_5_W0_en;
  wire  mem_60_5_W0_mask;
  wire [25:0] mem_60_6_R0_addr;
  wire  mem_60_6_R0_clk;
  wire [7:0] mem_60_6_R0_data;
  wire  mem_60_6_R0_en;
  wire [25:0] mem_60_6_W0_addr;
  wire  mem_60_6_W0_clk;
  wire [7:0] mem_60_6_W0_data;
  wire  mem_60_6_W0_en;
  wire  mem_60_6_W0_mask;
  wire [25:0] mem_60_7_R0_addr;
  wire  mem_60_7_R0_clk;
  wire [7:0] mem_60_7_R0_data;
  wire  mem_60_7_R0_en;
  wire [25:0] mem_60_7_W0_addr;
  wire  mem_60_7_W0_clk;
  wire [7:0] mem_60_7_W0_data;
  wire  mem_60_7_W0_en;
  wire  mem_60_7_W0_mask;
  wire [25:0] mem_61_0_R0_addr;
  wire  mem_61_0_R0_clk;
  wire [7:0] mem_61_0_R0_data;
  wire  mem_61_0_R0_en;
  wire [25:0] mem_61_0_W0_addr;
  wire  mem_61_0_W0_clk;
  wire [7:0] mem_61_0_W0_data;
  wire  mem_61_0_W0_en;
  wire  mem_61_0_W0_mask;
  wire [25:0] mem_61_1_R0_addr;
  wire  mem_61_1_R0_clk;
  wire [7:0] mem_61_1_R0_data;
  wire  mem_61_1_R0_en;
  wire [25:0] mem_61_1_W0_addr;
  wire  mem_61_1_W0_clk;
  wire [7:0] mem_61_1_W0_data;
  wire  mem_61_1_W0_en;
  wire  mem_61_1_W0_mask;
  wire [25:0] mem_61_2_R0_addr;
  wire  mem_61_2_R0_clk;
  wire [7:0] mem_61_2_R0_data;
  wire  mem_61_2_R0_en;
  wire [25:0] mem_61_2_W0_addr;
  wire  mem_61_2_W0_clk;
  wire [7:0] mem_61_2_W0_data;
  wire  mem_61_2_W0_en;
  wire  mem_61_2_W0_mask;
  wire [25:0] mem_61_3_R0_addr;
  wire  mem_61_3_R0_clk;
  wire [7:0] mem_61_3_R0_data;
  wire  mem_61_3_R0_en;
  wire [25:0] mem_61_3_W0_addr;
  wire  mem_61_3_W0_clk;
  wire [7:0] mem_61_3_W0_data;
  wire  mem_61_3_W0_en;
  wire  mem_61_3_W0_mask;
  wire [25:0] mem_61_4_R0_addr;
  wire  mem_61_4_R0_clk;
  wire [7:0] mem_61_4_R0_data;
  wire  mem_61_4_R0_en;
  wire [25:0] mem_61_4_W0_addr;
  wire  mem_61_4_W0_clk;
  wire [7:0] mem_61_4_W0_data;
  wire  mem_61_4_W0_en;
  wire  mem_61_4_W0_mask;
  wire [25:0] mem_61_5_R0_addr;
  wire  mem_61_5_R0_clk;
  wire [7:0] mem_61_5_R0_data;
  wire  mem_61_5_R0_en;
  wire [25:0] mem_61_5_W0_addr;
  wire  mem_61_5_W0_clk;
  wire [7:0] mem_61_5_W0_data;
  wire  mem_61_5_W0_en;
  wire  mem_61_5_W0_mask;
  wire [25:0] mem_61_6_R0_addr;
  wire  mem_61_6_R0_clk;
  wire [7:0] mem_61_6_R0_data;
  wire  mem_61_6_R0_en;
  wire [25:0] mem_61_6_W0_addr;
  wire  mem_61_6_W0_clk;
  wire [7:0] mem_61_6_W0_data;
  wire  mem_61_6_W0_en;
  wire  mem_61_6_W0_mask;
  wire [25:0] mem_61_7_R0_addr;
  wire  mem_61_7_R0_clk;
  wire [7:0] mem_61_7_R0_data;
  wire  mem_61_7_R0_en;
  wire [25:0] mem_61_7_W0_addr;
  wire  mem_61_7_W0_clk;
  wire [7:0] mem_61_7_W0_data;
  wire  mem_61_7_W0_en;
  wire  mem_61_7_W0_mask;
  wire [25:0] mem_62_0_R0_addr;
  wire  mem_62_0_R0_clk;
  wire [7:0] mem_62_0_R0_data;
  wire  mem_62_0_R0_en;
  wire [25:0] mem_62_0_W0_addr;
  wire  mem_62_0_W0_clk;
  wire [7:0] mem_62_0_W0_data;
  wire  mem_62_0_W0_en;
  wire  mem_62_0_W0_mask;
  wire [25:0] mem_62_1_R0_addr;
  wire  mem_62_1_R0_clk;
  wire [7:0] mem_62_1_R0_data;
  wire  mem_62_1_R0_en;
  wire [25:0] mem_62_1_W0_addr;
  wire  mem_62_1_W0_clk;
  wire [7:0] mem_62_1_W0_data;
  wire  mem_62_1_W0_en;
  wire  mem_62_1_W0_mask;
  wire [25:0] mem_62_2_R0_addr;
  wire  mem_62_2_R0_clk;
  wire [7:0] mem_62_2_R0_data;
  wire  mem_62_2_R0_en;
  wire [25:0] mem_62_2_W0_addr;
  wire  mem_62_2_W0_clk;
  wire [7:0] mem_62_2_W0_data;
  wire  mem_62_2_W0_en;
  wire  mem_62_2_W0_mask;
  wire [25:0] mem_62_3_R0_addr;
  wire  mem_62_3_R0_clk;
  wire [7:0] mem_62_3_R0_data;
  wire  mem_62_3_R0_en;
  wire [25:0] mem_62_3_W0_addr;
  wire  mem_62_3_W0_clk;
  wire [7:0] mem_62_3_W0_data;
  wire  mem_62_3_W0_en;
  wire  mem_62_3_W0_mask;
  wire [25:0] mem_62_4_R0_addr;
  wire  mem_62_4_R0_clk;
  wire [7:0] mem_62_4_R0_data;
  wire  mem_62_4_R0_en;
  wire [25:0] mem_62_4_W0_addr;
  wire  mem_62_4_W0_clk;
  wire [7:0] mem_62_4_W0_data;
  wire  mem_62_4_W0_en;
  wire  mem_62_4_W0_mask;
  wire [25:0] mem_62_5_R0_addr;
  wire  mem_62_5_R0_clk;
  wire [7:0] mem_62_5_R0_data;
  wire  mem_62_5_R0_en;
  wire [25:0] mem_62_5_W0_addr;
  wire  mem_62_5_W0_clk;
  wire [7:0] mem_62_5_W0_data;
  wire  mem_62_5_W0_en;
  wire  mem_62_5_W0_mask;
  wire [25:0] mem_62_6_R0_addr;
  wire  mem_62_6_R0_clk;
  wire [7:0] mem_62_6_R0_data;
  wire  mem_62_6_R0_en;
  wire [25:0] mem_62_6_W0_addr;
  wire  mem_62_6_W0_clk;
  wire [7:0] mem_62_6_W0_data;
  wire  mem_62_6_W0_en;
  wire  mem_62_6_W0_mask;
  wire [25:0] mem_62_7_R0_addr;
  wire  mem_62_7_R0_clk;
  wire [7:0] mem_62_7_R0_data;
  wire  mem_62_7_R0_en;
  wire [25:0] mem_62_7_W0_addr;
  wire  mem_62_7_W0_clk;
  wire [7:0] mem_62_7_W0_data;
  wire  mem_62_7_W0_en;
  wire  mem_62_7_W0_mask;
  wire [25:0] mem_63_0_R0_addr;
  wire  mem_63_0_R0_clk;
  wire [7:0] mem_63_0_R0_data;
  wire  mem_63_0_R0_en;
  wire [25:0] mem_63_0_W0_addr;
  wire  mem_63_0_W0_clk;
  wire [7:0] mem_63_0_W0_data;
  wire  mem_63_0_W0_en;
  wire  mem_63_0_W0_mask;
  wire [25:0] mem_63_1_R0_addr;
  wire  mem_63_1_R0_clk;
  wire [7:0] mem_63_1_R0_data;
  wire  mem_63_1_R0_en;
  wire [25:0] mem_63_1_W0_addr;
  wire  mem_63_1_W0_clk;
  wire [7:0] mem_63_1_W0_data;
  wire  mem_63_1_W0_en;
  wire  mem_63_1_W0_mask;
  wire [25:0] mem_63_2_R0_addr;
  wire  mem_63_2_R0_clk;
  wire [7:0] mem_63_2_R0_data;
  wire  mem_63_2_R0_en;
  wire [25:0] mem_63_2_W0_addr;
  wire  mem_63_2_W0_clk;
  wire [7:0] mem_63_2_W0_data;
  wire  mem_63_2_W0_en;
  wire  mem_63_2_W0_mask;
  wire [25:0] mem_63_3_R0_addr;
  wire  mem_63_3_R0_clk;
  wire [7:0] mem_63_3_R0_data;
  wire  mem_63_3_R0_en;
  wire [25:0] mem_63_3_W0_addr;
  wire  mem_63_3_W0_clk;
  wire [7:0] mem_63_3_W0_data;
  wire  mem_63_3_W0_en;
  wire  mem_63_3_W0_mask;
  wire [25:0] mem_63_4_R0_addr;
  wire  mem_63_4_R0_clk;
  wire [7:0] mem_63_4_R0_data;
  wire  mem_63_4_R0_en;
  wire [25:0] mem_63_4_W0_addr;
  wire  mem_63_4_W0_clk;
  wire [7:0] mem_63_4_W0_data;
  wire  mem_63_4_W0_en;
  wire  mem_63_4_W0_mask;
  wire [25:0] mem_63_5_R0_addr;
  wire  mem_63_5_R0_clk;
  wire [7:0] mem_63_5_R0_data;
  wire  mem_63_5_R0_en;
  wire [25:0] mem_63_5_W0_addr;
  wire  mem_63_5_W0_clk;
  wire [7:0] mem_63_5_W0_data;
  wire  mem_63_5_W0_en;
  wire  mem_63_5_W0_mask;
  wire [25:0] mem_63_6_R0_addr;
  wire  mem_63_6_R0_clk;
  wire [7:0] mem_63_6_R0_data;
  wire  mem_63_6_R0_en;
  wire [25:0] mem_63_6_W0_addr;
  wire  mem_63_6_W0_clk;
  wire [7:0] mem_63_6_W0_data;
  wire  mem_63_6_W0_en;
  wire  mem_63_6_W0_mask;
  wire [25:0] mem_63_7_R0_addr;
  wire  mem_63_7_R0_clk;
  wire [7:0] mem_63_7_R0_data;
  wire  mem_63_7_R0_en;
  wire [25:0] mem_63_7_W0_addr;
  wire  mem_63_7_W0_clk;
  wire [7:0] mem_63_7_W0_data;
  wire  mem_63_7_W0_en;
  wire  mem_63_7_W0_mask;
  wire [25:0] mem_64_0_R0_addr;
  wire  mem_64_0_R0_clk;
  wire [7:0] mem_64_0_R0_data;
  wire  mem_64_0_R0_en;
  wire [25:0] mem_64_0_W0_addr;
  wire  mem_64_0_W0_clk;
  wire [7:0] mem_64_0_W0_data;
  wire  mem_64_0_W0_en;
  wire  mem_64_0_W0_mask;
  wire [25:0] mem_64_1_R0_addr;
  wire  mem_64_1_R0_clk;
  wire [7:0] mem_64_1_R0_data;
  wire  mem_64_1_R0_en;
  wire [25:0] mem_64_1_W0_addr;
  wire  mem_64_1_W0_clk;
  wire [7:0] mem_64_1_W0_data;
  wire  mem_64_1_W0_en;
  wire  mem_64_1_W0_mask;
  wire [25:0] mem_64_2_R0_addr;
  wire  mem_64_2_R0_clk;
  wire [7:0] mem_64_2_R0_data;
  wire  mem_64_2_R0_en;
  wire [25:0] mem_64_2_W0_addr;
  wire  mem_64_2_W0_clk;
  wire [7:0] mem_64_2_W0_data;
  wire  mem_64_2_W0_en;
  wire  mem_64_2_W0_mask;
  wire [25:0] mem_64_3_R0_addr;
  wire  mem_64_3_R0_clk;
  wire [7:0] mem_64_3_R0_data;
  wire  mem_64_3_R0_en;
  wire [25:0] mem_64_3_W0_addr;
  wire  mem_64_3_W0_clk;
  wire [7:0] mem_64_3_W0_data;
  wire  mem_64_3_W0_en;
  wire  mem_64_3_W0_mask;
  wire [25:0] mem_64_4_R0_addr;
  wire  mem_64_4_R0_clk;
  wire [7:0] mem_64_4_R0_data;
  wire  mem_64_4_R0_en;
  wire [25:0] mem_64_4_W0_addr;
  wire  mem_64_4_W0_clk;
  wire [7:0] mem_64_4_W0_data;
  wire  mem_64_4_W0_en;
  wire  mem_64_4_W0_mask;
  wire [25:0] mem_64_5_R0_addr;
  wire  mem_64_5_R0_clk;
  wire [7:0] mem_64_5_R0_data;
  wire  mem_64_5_R0_en;
  wire [25:0] mem_64_5_W0_addr;
  wire  mem_64_5_W0_clk;
  wire [7:0] mem_64_5_W0_data;
  wire  mem_64_5_W0_en;
  wire  mem_64_5_W0_mask;
  wire [25:0] mem_64_6_R0_addr;
  wire  mem_64_6_R0_clk;
  wire [7:0] mem_64_6_R0_data;
  wire  mem_64_6_R0_en;
  wire [25:0] mem_64_6_W0_addr;
  wire  mem_64_6_W0_clk;
  wire [7:0] mem_64_6_W0_data;
  wire  mem_64_6_W0_en;
  wire  mem_64_6_W0_mask;
  wire [25:0] mem_64_7_R0_addr;
  wire  mem_64_7_R0_clk;
  wire [7:0] mem_64_7_R0_data;
  wire  mem_64_7_R0_en;
  wire [25:0] mem_64_7_W0_addr;
  wire  mem_64_7_W0_clk;
  wire [7:0] mem_64_7_W0_data;
  wire  mem_64_7_W0_en;
  wire  mem_64_7_W0_mask;
  wire [25:0] mem_65_0_R0_addr;
  wire  mem_65_0_R0_clk;
  wire [7:0] mem_65_0_R0_data;
  wire  mem_65_0_R0_en;
  wire [25:0] mem_65_0_W0_addr;
  wire  mem_65_0_W0_clk;
  wire [7:0] mem_65_0_W0_data;
  wire  mem_65_0_W0_en;
  wire  mem_65_0_W0_mask;
  wire [25:0] mem_65_1_R0_addr;
  wire  mem_65_1_R0_clk;
  wire [7:0] mem_65_1_R0_data;
  wire  mem_65_1_R0_en;
  wire [25:0] mem_65_1_W0_addr;
  wire  mem_65_1_W0_clk;
  wire [7:0] mem_65_1_W0_data;
  wire  mem_65_1_W0_en;
  wire  mem_65_1_W0_mask;
  wire [25:0] mem_65_2_R0_addr;
  wire  mem_65_2_R0_clk;
  wire [7:0] mem_65_2_R0_data;
  wire  mem_65_2_R0_en;
  wire [25:0] mem_65_2_W0_addr;
  wire  mem_65_2_W0_clk;
  wire [7:0] mem_65_2_W0_data;
  wire  mem_65_2_W0_en;
  wire  mem_65_2_W0_mask;
  wire [25:0] mem_65_3_R0_addr;
  wire  mem_65_3_R0_clk;
  wire [7:0] mem_65_3_R0_data;
  wire  mem_65_3_R0_en;
  wire [25:0] mem_65_3_W0_addr;
  wire  mem_65_3_W0_clk;
  wire [7:0] mem_65_3_W0_data;
  wire  mem_65_3_W0_en;
  wire  mem_65_3_W0_mask;
  wire [25:0] mem_65_4_R0_addr;
  wire  mem_65_4_R0_clk;
  wire [7:0] mem_65_4_R0_data;
  wire  mem_65_4_R0_en;
  wire [25:0] mem_65_4_W0_addr;
  wire  mem_65_4_W0_clk;
  wire [7:0] mem_65_4_W0_data;
  wire  mem_65_4_W0_en;
  wire  mem_65_4_W0_mask;
  wire [25:0] mem_65_5_R0_addr;
  wire  mem_65_5_R0_clk;
  wire [7:0] mem_65_5_R0_data;
  wire  mem_65_5_R0_en;
  wire [25:0] mem_65_5_W0_addr;
  wire  mem_65_5_W0_clk;
  wire [7:0] mem_65_5_W0_data;
  wire  mem_65_5_W0_en;
  wire  mem_65_5_W0_mask;
  wire [25:0] mem_65_6_R0_addr;
  wire  mem_65_6_R0_clk;
  wire [7:0] mem_65_6_R0_data;
  wire  mem_65_6_R0_en;
  wire [25:0] mem_65_6_W0_addr;
  wire  mem_65_6_W0_clk;
  wire [7:0] mem_65_6_W0_data;
  wire  mem_65_6_W0_en;
  wire  mem_65_6_W0_mask;
  wire [25:0] mem_65_7_R0_addr;
  wire  mem_65_7_R0_clk;
  wire [7:0] mem_65_7_R0_data;
  wire  mem_65_7_R0_en;
  wire [25:0] mem_65_7_W0_addr;
  wire  mem_65_7_W0_clk;
  wire [7:0] mem_65_7_W0_data;
  wire  mem_65_7_W0_en;
  wire  mem_65_7_W0_mask;
  wire [25:0] mem_66_0_R0_addr;
  wire  mem_66_0_R0_clk;
  wire [7:0] mem_66_0_R0_data;
  wire  mem_66_0_R0_en;
  wire [25:0] mem_66_0_W0_addr;
  wire  mem_66_0_W0_clk;
  wire [7:0] mem_66_0_W0_data;
  wire  mem_66_0_W0_en;
  wire  mem_66_0_W0_mask;
  wire [25:0] mem_66_1_R0_addr;
  wire  mem_66_1_R0_clk;
  wire [7:0] mem_66_1_R0_data;
  wire  mem_66_1_R0_en;
  wire [25:0] mem_66_1_W0_addr;
  wire  mem_66_1_W0_clk;
  wire [7:0] mem_66_1_W0_data;
  wire  mem_66_1_W0_en;
  wire  mem_66_1_W0_mask;
  wire [25:0] mem_66_2_R0_addr;
  wire  mem_66_2_R0_clk;
  wire [7:0] mem_66_2_R0_data;
  wire  mem_66_2_R0_en;
  wire [25:0] mem_66_2_W0_addr;
  wire  mem_66_2_W0_clk;
  wire [7:0] mem_66_2_W0_data;
  wire  mem_66_2_W0_en;
  wire  mem_66_2_W0_mask;
  wire [25:0] mem_66_3_R0_addr;
  wire  mem_66_3_R0_clk;
  wire [7:0] mem_66_3_R0_data;
  wire  mem_66_3_R0_en;
  wire [25:0] mem_66_3_W0_addr;
  wire  mem_66_3_W0_clk;
  wire [7:0] mem_66_3_W0_data;
  wire  mem_66_3_W0_en;
  wire  mem_66_3_W0_mask;
  wire [25:0] mem_66_4_R0_addr;
  wire  mem_66_4_R0_clk;
  wire [7:0] mem_66_4_R0_data;
  wire  mem_66_4_R0_en;
  wire [25:0] mem_66_4_W0_addr;
  wire  mem_66_4_W0_clk;
  wire [7:0] mem_66_4_W0_data;
  wire  mem_66_4_W0_en;
  wire  mem_66_4_W0_mask;
  wire [25:0] mem_66_5_R0_addr;
  wire  mem_66_5_R0_clk;
  wire [7:0] mem_66_5_R0_data;
  wire  mem_66_5_R0_en;
  wire [25:0] mem_66_5_W0_addr;
  wire  mem_66_5_W0_clk;
  wire [7:0] mem_66_5_W0_data;
  wire  mem_66_5_W0_en;
  wire  mem_66_5_W0_mask;
  wire [25:0] mem_66_6_R0_addr;
  wire  mem_66_6_R0_clk;
  wire [7:0] mem_66_6_R0_data;
  wire  mem_66_6_R0_en;
  wire [25:0] mem_66_6_W0_addr;
  wire  mem_66_6_W0_clk;
  wire [7:0] mem_66_6_W0_data;
  wire  mem_66_6_W0_en;
  wire  mem_66_6_W0_mask;
  wire [25:0] mem_66_7_R0_addr;
  wire  mem_66_7_R0_clk;
  wire [7:0] mem_66_7_R0_data;
  wire  mem_66_7_R0_en;
  wire [25:0] mem_66_7_W0_addr;
  wire  mem_66_7_W0_clk;
  wire [7:0] mem_66_7_W0_data;
  wire  mem_66_7_W0_en;
  wire  mem_66_7_W0_mask;
  wire [25:0] mem_67_0_R0_addr;
  wire  mem_67_0_R0_clk;
  wire [7:0] mem_67_0_R0_data;
  wire  mem_67_0_R0_en;
  wire [25:0] mem_67_0_W0_addr;
  wire  mem_67_0_W0_clk;
  wire [7:0] mem_67_0_W0_data;
  wire  mem_67_0_W0_en;
  wire  mem_67_0_W0_mask;
  wire [25:0] mem_67_1_R0_addr;
  wire  mem_67_1_R0_clk;
  wire [7:0] mem_67_1_R0_data;
  wire  mem_67_1_R0_en;
  wire [25:0] mem_67_1_W0_addr;
  wire  mem_67_1_W0_clk;
  wire [7:0] mem_67_1_W0_data;
  wire  mem_67_1_W0_en;
  wire  mem_67_1_W0_mask;
  wire [25:0] mem_67_2_R0_addr;
  wire  mem_67_2_R0_clk;
  wire [7:0] mem_67_2_R0_data;
  wire  mem_67_2_R0_en;
  wire [25:0] mem_67_2_W0_addr;
  wire  mem_67_2_W0_clk;
  wire [7:0] mem_67_2_W0_data;
  wire  mem_67_2_W0_en;
  wire  mem_67_2_W0_mask;
  wire [25:0] mem_67_3_R0_addr;
  wire  mem_67_3_R0_clk;
  wire [7:0] mem_67_3_R0_data;
  wire  mem_67_3_R0_en;
  wire [25:0] mem_67_3_W0_addr;
  wire  mem_67_3_W0_clk;
  wire [7:0] mem_67_3_W0_data;
  wire  mem_67_3_W0_en;
  wire  mem_67_3_W0_mask;
  wire [25:0] mem_67_4_R0_addr;
  wire  mem_67_4_R0_clk;
  wire [7:0] mem_67_4_R0_data;
  wire  mem_67_4_R0_en;
  wire [25:0] mem_67_4_W0_addr;
  wire  mem_67_4_W0_clk;
  wire [7:0] mem_67_4_W0_data;
  wire  mem_67_4_W0_en;
  wire  mem_67_4_W0_mask;
  wire [25:0] mem_67_5_R0_addr;
  wire  mem_67_5_R0_clk;
  wire [7:0] mem_67_5_R0_data;
  wire  mem_67_5_R0_en;
  wire [25:0] mem_67_5_W0_addr;
  wire  mem_67_5_W0_clk;
  wire [7:0] mem_67_5_W0_data;
  wire  mem_67_5_W0_en;
  wire  mem_67_5_W0_mask;
  wire [25:0] mem_67_6_R0_addr;
  wire  mem_67_6_R0_clk;
  wire [7:0] mem_67_6_R0_data;
  wire  mem_67_6_R0_en;
  wire [25:0] mem_67_6_W0_addr;
  wire  mem_67_6_W0_clk;
  wire [7:0] mem_67_6_W0_data;
  wire  mem_67_6_W0_en;
  wire  mem_67_6_W0_mask;
  wire [25:0] mem_67_7_R0_addr;
  wire  mem_67_7_R0_clk;
  wire [7:0] mem_67_7_R0_data;
  wire  mem_67_7_R0_en;
  wire [25:0] mem_67_7_W0_addr;
  wire  mem_67_7_W0_clk;
  wire [7:0] mem_67_7_W0_data;
  wire  mem_67_7_W0_en;
  wire  mem_67_7_W0_mask;
  wire [25:0] mem_68_0_R0_addr;
  wire  mem_68_0_R0_clk;
  wire [7:0] mem_68_0_R0_data;
  wire  mem_68_0_R0_en;
  wire [25:0] mem_68_0_W0_addr;
  wire  mem_68_0_W0_clk;
  wire [7:0] mem_68_0_W0_data;
  wire  mem_68_0_W0_en;
  wire  mem_68_0_W0_mask;
  wire [25:0] mem_68_1_R0_addr;
  wire  mem_68_1_R0_clk;
  wire [7:0] mem_68_1_R0_data;
  wire  mem_68_1_R0_en;
  wire [25:0] mem_68_1_W0_addr;
  wire  mem_68_1_W0_clk;
  wire [7:0] mem_68_1_W0_data;
  wire  mem_68_1_W0_en;
  wire  mem_68_1_W0_mask;
  wire [25:0] mem_68_2_R0_addr;
  wire  mem_68_2_R0_clk;
  wire [7:0] mem_68_2_R0_data;
  wire  mem_68_2_R0_en;
  wire [25:0] mem_68_2_W0_addr;
  wire  mem_68_2_W0_clk;
  wire [7:0] mem_68_2_W0_data;
  wire  mem_68_2_W0_en;
  wire  mem_68_2_W0_mask;
  wire [25:0] mem_68_3_R0_addr;
  wire  mem_68_3_R0_clk;
  wire [7:0] mem_68_3_R0_data;
  wire  mem_68_3_R0_en;
  wire [25:0] mem_68_3_W0_addr;
  wire  mem_68_3_W0_clk;
  wire [7:0] mem_68_3_W0_data;
  wire  mem_68_3_W0_en;
  wire  mem_68_3_W0_mask;
  wire [25:0] mem_68_4_R0_addr;
  wire  mem_68_4_R0_clk;
  wire [7:0] mem_68_4_R0_data;
  wire  mem_68_4_R0_en;
  wire [25:0] mem_68_4_W0_addr;
  wire  mem_68_4_W0_clk;
  wire [7:0] mem_68_4_W0_data;
  wire  mem_68_4_W0_en;
  wire  mem_68_4_W0_mask;
  wire [25:0] mem_68_5_R0_addr;
  wire  mem_68_5_R0_clk;
  wire [7:0] mem_68_5_R0_data;
  wire  mem_68_5_R0_en;
  wire [25:0] mem_68_5_W0_addr;
  wire  mem_68_5_W0_clk;
  wire [7:0] mem_68_5_W0_data;
  wire  mem_68_5_W0_en;
  wire  mem_68_5_W0_mask;
  wire [25:0] mem_68_6_R0_addr;
  wire  mem_68_6_R0_clk;
  wire [7:0] mem_68_6_R0_data;
  wire  mem_68_6_R0_en;
  wire [25:0] mem_68_6_W0_addr;
  wire  mem_68_6_W0_clk;
  wire [7:0] mem_68_6_W0_data;
  wire  mem_68_6_W0_en;
  wire  mem_68_6_W0_mask;
  wire [25:0] mem_68_7_R0_addr;
  wire  mem_68_7_R0_clk;
  wire [7:0] mem_68_7_R0_data;
  wire  mem_68_7_R0_en;
  wire [25:0] mem_68_7_W0_addr;
  wire  mem_68_7_W0_clk;
  wire [7:0] mem_68_7_W0_data;
  wire  mem_68_7_W0_en;
  wire  mem_68_7_W0_mask;
  wire [25:0] mem_69_0_R0_addr;
  wire  mem_69_0_R0_clk;
  wire [7:0] mem_69_0_R0_data;
  wire  mem_69_0_R0_en;
  wire [25:0] mem_69_0_W0_addr;
  wire  mem_69_0_W0_clk;
  wire [7:0] mem_69_0_W0_data;
  wire  mem_69_0_W0_en;
  wire  mem_69_0_W0_mask;
  wire [25:0] mem_69_1_R0_addr;
  wire  mem_69_1_R0_clk;
  wire [7:0] mem_69_1_R0_data;
  wire  mem_69_1_R0_en;
  wire [25:0] mem_69_1_W0_addr;
  wire  mem_69_1_W0_clk;
  wire [7:0] mem_69_1_W0_data;
  wire  mem_69_1_W0_en;
  wire  mem_69_1_W0_mask;
  wire [25:0] mem_69_2_R0_addr;
  wire  mem_69_2_R0_clk;
  wire [7:0] mem_69_2_R0_data;
  wire  mem_69_2_R0_en;
  wire [25:0] mem_69_2_W0_addr;
  wire  mem_69_2_W0_clk;
  wire [7:0] mem_69_2_W0_data;
  wire  mem_69_2_W0_en;
  wire  mem_69_2_W0_mask;
  wire [25:0] mem_69_3_R0_addr;
  wire  mem_69_3_R0_clk;
  wire [7:0] mem_69_3_R0_data;
  wire  mem_69_3_R0_en;
  wire [25:0] mem_69_3_W0_addr;
  wire  mem_69_3_W0_clk;
  wire [7:0] mem_69_3_W0_data;
  wire  mem_69_3_W0_en;
  wire  mem_69_3_W0_mask;
  wire [25:0] mem_69_4_R0_addr;
  wire  mem_69_4_R0_clk;
  wire [7:0] mem_69_4_R0_data;
  wire  mem_69_4_R0_en;
  wire [25:0] mem_69_4_W0_addr;
  wire  mem_69_4_W0_clk;
  wire [7:0] mem_69_4_W0_data;
  wire  mem_69_4_W0_en;
  wire  mem_69_4_W0_mask;
  wire [25:0] mem_69_5_R0_addr;
  wire  mem_69_5_R0_clk;
  wire [7:0] mem_69_5_R0_data;
  wire  mem_69_5_R0_en;
  wire [25:0] mem_69_5_W0_addr;
  wire  mem_69_5_W0_clk;
  wire [7:0] mem_69_5_W0_data;
  wire  mem_69_5_W0_en;
  wire  mem_69_5_W0_mask;
  wire [25:0] mem_69_6_R0_addr;
  wire  mem_69_6_R0_clk;
  wire [7:0] mem_69_6_R0_data;
  wire  mem_69_6_R0_en;
  wire [25:0] mem_69_6_W0_addr;
  wire  mem_69_6_W0_clk;
  wire [7:0] mem_69_6_W0_data;
  wire  mem_69_6_W0_en;
  wire  mem_69_6_W0_mask;
  wire [25:0] mem_69_7_R0_addr;
  wire  mem_69_7_R0_clk;
  wire [7:0] mem_69_7_R0_data;
  wire  mem_69_7_R0_en;
  wire [25:0] mem_69_7_W0_addr;
  wire  mem_69_7_W0_clk;
  wire [7:0] mem_69_7_W0_data;
  wire  mem_69_7_W0_en;
  wire  mem_69_7_W0_mask;
  wire [25:0] mem_70_0_R0_addr;
  wire  mem_70_0_R0_clk;
  wire [7:0] mem_70_0_R0_data;
  wire  mem_70_0_R0_en;
  wire [25:0] mem_70_0_W0_addr;
  wire  mem_70_0_W0_clk;
  wire [7:0] mem_70_0_W0_data;
  wire  mem_70_0_W0_en;
  wire  mem_70_0_W0_mask;
  wire [25:0] mem_70_1_R0_addr;
  wire  mem_70_1_R0_clk;
  wire [7:0] mem_70_1_R0_data;
  wire  mem_70_1_R0_en;
  wire [25:0] mem_70_1_W0_addr;
  wire  mem_70_1_W0_clk;
  wire [7:0] mem_70_1_W0_data;
  wire  mem_70_1_W0_en;
  wire  mem_70_1_W0_mask;
  wire [25:0] mem_70_2_R0_addr;
  wire  mem_70_2_R0_clk;
  wire [7:0] mem_70_2_R0_data;
  wire  mem_70_2_R0_en;
  wire [25:0] mem_70_2_W0_addr;
  wire  mem_70_2_W0_clk;
  wire [7:0] mem_70_2_W0_data;
  wire  mem_70_2_W0_en;
  wire  mem_70_2_W0_mask;
  wire [25:0] mem_70_3_R0_addr;
  wire  mem_70_3_R0_clk;
  wire [7:0] mem_70_3_R0_data;
  wire  mem_70_3_R0_en;
  wire [25:0] mem_70_3_W0_addr;
  wire  mem_70_3_W0_clk;
  wire [7:0] mem_70_3_W0_data;
  wire  mem_70_3_W0_en;
  wire  mem_70_3_W0_mask;
  wire [25:0] mem_70_4_R0_addr;
  wire  mem_70_4_R0_clk;
  wire [7:0] mem_70_4_R0_data;
  wire  mem_70_4_R0_en;
  wire [25:0] mem_70_4_W0_addr;
  wire  mem_70_4_W0_clk;
  wire [7:0] mem_70_4_W0_data;
  wire  mem_70_4_W0_en;
  wire  mem_70_4_W0_mask;
  wire [25:0] mem_70_5_R0_addr;
  wire  mem_70_5_R0_clk;
  wire [7:0] mem_70_5_R0_data;
  wire  mem_70_5_R0_en;
  wire [25:0] mem_70_5_W0_addr;
  wire  mem_70_5_W0_clk;
  wire [7:0] mem_70_5_W0_data;
  wire  mem_70_5_W0_en;
  wire  mem_70_5_W0_mask;
  wire [25:0] mem_70_6_R0_addr;
  wire  mem_70_6_R0_clk;
  wire [7:0] mem_70_6_R0_data;
  wire  mem_70_6_R0_en;
  wire [25:0] mem_70_6_W0_addr;
  wire  mem_70_6_W0_clk;
  wire [7:0] mem_70_6_W0_data;
  wire  mem_70_6_W0_en;
  wire  mem_70_6_W0_mask;
  wire [25:0] mem_70_7_R0_addr;
  wire  mem_70_7_R0_clk;
  wire [7:0] mem_70_7_R0_data;
  wire  mem_70_7_R0_en;
  wire [25:0] mem_70_7_W0_addr;
  wire  mem_70_7_W0_clk;
  wire [7:0] mem_70_7_W0_data;
  wire  mem_70_7_W0_en;
  wire  mem_70_7_W0_mask;
  wire [25:0] mem_71_0_R0_addr;
  wire  mem_71_0_R0_clk;
  wire [7:0] mem_71_0_R0_data;
  wire  mem_71_0_R0_en;
  wire [25:0] mem_71_0_W0_addr;
  wire  mem_71_0_W0_clk;
  wire [7:0] mem_71_0_W0_data;
  wire  mem_71_0_W0_en;
  wire  mem_71_0_W0_mask;
  wire [25:0] mem_71_1_R0_addr;
  wire  mem_71_1_R0_clk;
  wire [7:0] mem_71_1_R0_data;
  wire  mem_71_1_R0_en;
  wire [25:0] mem_71_1_W0_addr;
  wire  mem_71_1_W0_clk;
  wire [7:0] mem_71_1_W0_data;
  wire  mem_71_1_W0_en;
  wire  mem_71_1_W0_mask;
  wire [25:0] mem_71_2_R0_addr;
  wire  mem_71_2_R0_clk;
  wire [7:0] mem_71_2_R0_data;
  wire  mem_71_2_R0_en;
  wire [25:0] mem_71_2_W0_addr;
  wire  mem_71_2_W0_clk;
  wire [7:0] mem_71_2_W0_data;
  wire  mem_71_2_W0_en;
  wire  mem_71_2_W0_mask;
  wire [25:0] mem_71_3_R0_addr;
  wire  mem_71_3_R0_clk;
  wire [7:0] mem_71_3_R0_data;
  wire  mem_71_3_R0_en;
  wire [25:0] mem_71_3_W0_addr;
  wire  mem_71_3_W0_clk;
  wire [7:0] mem_71_3_W0_data;
  wire  mem_71_3_W0_en;
  wire  mem_71_3_W0_mask;
  wire [25:0] mem_71_4_R0_addr;
  wire  mem_71_4_R0_clk;
  wire [7:0] mem_71_4_R0_data;
  wire  mem_71_4_R0_en;
  wire [25:0] mem_71_4_W0_addr;
  wire  mem_71_4_W0_clk;
  wire [7:0] mem_71_4_W0_data;
  wire  mem_71_4_W0_en;
  wire  mem_71_4_W0_mask;
  wire [25:0] mem_71_5_R0_addr;
  wire  mem_71_5_R0_clk;
  wire [7:0] mem_71_5_R0_data;
  wire  mem_71_5_R0_en;
  wire [25:0] mem_71_5_W0_addr;
  wire  mem_71_5_W0_clk;
  wire [7:0] mem_71_5_W0_data;
  wire  mem_71_5_W0_en;
  wire  mem_71_5_W0_mask;
  wire [25:0] mem_71_6_R0_addr;
  wire  mem_71_6_R0_clk;
  wire [7:0] mem_71_6_R0_data;
  wire  mem_71_6_R0_en;
  wire [25:0] mem_71_6_W0_addr;
  wire  mem_71_6_W0_clk;
  wire [7:0] mem_71_6_W0_data;
  wire  mem_71_6_W0_en;
  wire  mem_71_6_W0_mask;
  wire [25:0] mem_71_7_R0_addr;
  wire  mem_71_7_R0_clk;
  wire [7:0] mem_71_7_R0_data;
  wire  mem_71_7_R0_en;
  wire [25:0] mem_71_7_W0_addr;
  wire  mem_71_7_W0_clk;
  wire [7:0] mem_71_7_W0_data;
  wire  mem_71_7_W0_en;
  wire  mem_71_7_W0_mask;
  wire [25:0] mem_72_0_R0_addr;
  wire  mem_72_0_R0_clk;
  wire [7:0] mem_72_0_R0_data;
  wire  mem_72_0_R0_en;
  wire [25:0] mem_72_0_W0_addr;
  wire  mem_72_0_W0_clk;
  wire [7:0] mem_72_0_W0_data;
  wire  mem_72_0_W0_en;
  wire  mem_72_0_W0_mask;
  wire [25:0] mem_72_1_R0_addr;
  wire  mem_72_1_R0_clk;
  wire [7:0] mem_72_1_R0_data;
  wire  mem_72_1_R0_en;
  wire [25:0] mem_72_1_W0_addr;
  wire  mem_72_1_W0_clk;
  wire [7:0] mem_72_1_W0_data;
  wire  mem_72_1_W0_en;
  wire  mem_72_1_W0_mask;
  wire [25:0] mem_72_2_R0_addr;
  wire  mem_72_2_R0_clk;
  wire [7:0] mem_72_2_R0_data;
  wire  mem_72_2_R0_en;
  wire [25:0] mem_72_2_W0_addr;
  wire  mem_72_2_W0_clk;
  wire [7:0] mem_72_2_W0_data;
  wire  mem_72_2_W0_en;
  wire  mem_72_2_W0_mask;
  wire [25:0] mem_72_3_R0_addr;
  wire  mem_72_3_R0_clk;
  wire [7:0] mem_72_3_R0_data;
  wire  mem_72_3_R0_en;
  wire [25:0] mem_72_3_W0_addr;
  wire  mem_72_3_W0_clk;
  wire [7:0] mem_72_3_W0_data;
  wire  mem_72_3_W0_en;
  wire  mem_72_3_W0_mask;
  wire [25:0] mem_72_4_R0_addr;
  wire  mem_72_4_R0_clk;
  wire [7:0] mem_72_4_R0_data;
  wire  mem_72_4_R0_en;
  wire [25:0] mem_72_4_W0_addr;
  wire  mem_72_4_W0_clk;
  wire [7:0] mem_72_4_W0_data;
  wire  mem_72_4_W0_en;
  wire  mem_72_4_W0_mask;
  wire [25:0] mem_72_5_R0_addr;
  wire  mem_72_5_R0_clk;
  wire [7:0] mem_72_5_R0_data;
  wire  mem_72_5_R0_en;
  wire [25:0] mem_72_5_W0_addr;
  wire  mem_72_5_W0_clk;
  wire [7:0] mem_72_5_W0_data;
  wire  mem_72_5_W0_en;
  wire  mem_72_5_W0_mask;
  wire [25:0] mem_72_6_R0_addr;
  wire  mem_72_6_R0_clk;
  wire [7:0] mem_72_6_R0_data;
  wire  mem_72_6_R0_en;
  wire [25:0] mem_72_6_W0_addr;
  wire  mem_72_6_W0_clk;
  wire [7:0] mem_72_6_W0_data;
  wire  mem_72_6_W0_en;
  wire  mem_72_6_W0_mask;
  wire [25:0] mem_72_7_R0_addr;
  wire  mem_72_7_R0_clk;
  wire [7:0] mem_72_7_R0_data;
  wire  mem_72_7_R0_en;
  wire [25:0] mem_72_7_W0_addr;
  wire  mem_72_7_W0_clk;
  wire [7:0] mem_72_7_W0_data;
  wire  mem_72_7_W0_en;
  wire  mem_72_7_W0_mask;
  wire [25:0] mem_73_0_R0_addr;
  wire  mem_73_0_R0_clk;
  wire [7:0] mem_73_0_R0_data;
  wire  mem_73_0_R0_en;
  wire [25:0] mem_73_0_W0_addr;
  wire  mem_73_0_W0_clk;
  wire [7:0] mem_73_0_W0_data;
  wire  mem_73_0_W0_en;
  wire  mem_73_0_W0_mask;
  wire [25:0] mem_73_1_R0_addr;
  wire  mem_73_1_R0_clk;
  wire [7:0] mem_73_1_R0_data;
  wire  mem_73_1_R0_en;
  wire [25:0] mem_73_1_W0_addr;
  wire  mem_73_1_W0_clk;
  wire [7:0] mem_73_1_W0_data;
  wire  mem_73_1_W0_en;
  wire  mem_73_1_W0_mask;
  wire [25:0] mem_73_2_R0_addr;
  wire  mem_73_2_R0_clk;
  wire [7:0] mem_73_2_R0_data;
  wire  mem_73_2_R0_en;
  wire [25:0] mem_73_2_W0_addr;
  wire  mem_73_2_W0_clk;
  wire [7:0] mem_73_2_W0_data;
  wire  mem_73_2_W0_en;
  wire  mem_73_2_W0_mask;
  wire [25:0] mem_73_3_R0_addr;
  wire  mem_73_3_R0_clk;
  wire [7:0] mem_73_3_R0_data;
  wire  mem_73_3_R0_en;
  wire [25:0] mem_73_3_W0_addr;
  wire  mem_73_3_W0_clk;
  wire [7:0] mem_73_3_W0_data;
  wire  mem_73_3_W0_en;
  wire  mem_73_3_W0_mask;
  wire [25:0] mem_73_4_R0_addr;
  wire  mem_73_4_R0_clk;
  wire [7:0] mem_73_4_R0_data;
  wire  mem_73_4_R0_en;
  wire [25:0] mem_73_4_W0_addr;
  wire  mem_73_4_W0_clk;
  wire [7:0] mem_73_4_W0_data;
  wire  mem_73_4_W0_en;
  wire  mem_73_4_W0_mask;
  wire [25:0] mem_73_5_R0_addr;
  wire  mem_73_5_R0_clk;
  wire [7:0] mem_73_5_R0_data;
  wire  mem_73_5_R0_en;
  wire [25:0] mem_73_5_W0_addr;
  wire  mem_73_5_W0_clk;
  wire [7:0] mem_73_5_W0_data;
  wire  mem_73_5_W0_en;
  wire  mem_73_5_W0_mask;
  wire [25:0] mem_73_6_R0_addr;
  wire  mem_73_6_R0_clk;
  wire [7:0] mem_73_6_R0_data;
  wire  mem_73_6_R0_en;
  wire [25:0] mem_73_6_W0_addr;
  wire  mem_73_6_W0_clk;
  wire [7:0] mem_73_6_W0_data;
  wire  mem_73_6_W0_en;
  wire  mem_73_6_W0_mask;
  wire [25:0] mem_73_7_R0_addr;
  wire  mem_73_7_R0_clk;
  wire [7:0] mem_73_7_R0_data;
  wire  mem_73_7_R0_en;
  wire [25:0] mem_73_7_W0_addr;
  wire  mem_73_7_W0_clk;
  wire [7:0] mem_73_7_W0_data;
  wire  mem_73_7_W0_en;
  wire  mem_73_7_W0_mask;
  wire [25:0] mem_74_0_R0_addr;
  wire  mem_74_0_R0_clk;
  wire [7:0] mem_74_0_R0_data;
  wire  mem_74_0_R0_en;
  wire [25:0] mem_74_0_W0_addr;
  wire  mem_74_0_W0_clk;
  wire [7:0] mem_74_0_W0_data;
  wire  mem_74_0_W0_en;
  wire  mem_74_0_W0_mask;
  wire [25:0] mem_74_1_R0_addr;
  wire  mem_74_1_R0_clk;
  wire [7:0] mem_74_1_R0_data;
  wire  mem_74_1_R0_en;
  wire [25:0] mem_74_1_W0_addr;
  wire  mem_74_1_W0_clk;
  wire [7:0] mem_74_1_W0_data;
  wire  mem_74_1_W0_en;
  wire  mem_74_1_W0_mask;
  wire [25:0] mem_74_2_R0_addr;
  wire  mem_74_2_R0_clk;
  wire [7:0] mem_74_2_R0_data;
  wire  mem_74_2_R0_en;
  wire [25:0] mem_74_2_W0_addr;
  wire  mem_74_2_W0_clk;
  wire [7:0] mem_74_2_W0_data;
  wire  mem_74_2_W0_en;
  wire  mem_74_2_W0_mask;
  wire [25:0] mem_74_3_R0_addr;
  wire  mem_74_3_R0_clk;
  wire [7:0] mem_74_3_R0_data;
  wire  mem_74_3_R0_en;
  wire [25:0] mem_74_3_W0_addr;
  wire  mem_74_3_W0_clk;
  wire [7:0] mem_74_3_W0_data;
  wire  mem_74_3_W0_en;
  wire  mem_74_3_W0_mask;
  wire [25:0] mem_74_4_R0_addr;
  wire  mem_74_4_R0_clk;
  wire [7:0] mem_74_4_R0_data;
  wire  mem_74_4_R0_en;
  wire [25:0] mem_74_4_W0_addr;
  wire  mem_74_4_W0_clk;
  wire [7:0] mem_74_4_W0_data;
  wire  mem_74_4_W0_en;
  wire  mem_74_4_W0_mask;
  wire [25:0] mem_74_5_R0_addr;
  wire  mem_74_5_R0_clk;
  wire [7:0] mem_74_5_R0_data;
  wire  mem_74_5_R0_en;
  wire [25:0] mem_74_5_W0_addr;
  wire  mem_74_5_W0_clk;
  wire [7:0] mem_74_5_W0_data;
  wire  mem_74_5_W0_en;
  wire  mem_74_5_W0_mask;
  wire [25:0] mem_74_6_R0_addr;
  wire  mem_74_6_R0_clk;
  wire [7:0] mem_74_6_R0_data;
  wire  mem_74_6_R0_en;
  wire [25:0] mem_74_6_W0_addr;
  wire  mem_74_6_W0_clk;
  wire [7:0] mem_74_6_W0_data;
  wire  mem_74_6_W0_en;
  wire  mem_74_6_W0_mask;
  wire [25:0] mem_74_7_R0_addr;
  wire  mem_74_7_R0_clk;
  wire [7:0] mem_74_7_R0_data;
  wire  mem_74_7_R0_en;
  wire [25:0] mem_74_7_W0_addr;
  wire  mem_74_7_W0_clk;
  wire [7:0] mem_74_7_W0_data;
  wire  mem_74_7_W0_en;
  wire  mem_74_7_W0_mask;
  wire [25:0] mem_75_0_R0_addr;
  wire  mem_75_0_R0_clk;
  wire [7:0] mem_75_0_R0_data;
  wire  mem_75_0_R0_en;
  wire [25:0] mem_75_0_W0_addr;
  wire  mem_75_0_W0_clk;
  wire [7:0] mem_75_0_W0_data;
  wire  mem_75_0_W0_en;
  wire  mem_75_0_W0_mask;
  wire [25:0] mem_75_1_R0_addr;
  wire  mem_75_1_R0_clk;
  wire [7:0] mem_75_1_R0_data;
  wire  mem_75_1_R0_en;
  wire [25:0] mem_75_1_W0_addr;
  wire  mem_75_1_W0_clk;
  wire [7:0] mem_75_1_W0_data;
  wire  mem_75_1_W0_en;
  wire  mem_75_1_W0_mask;
  wire [25:0] mem_75_2_R0_addr;
  wire  mem_75_2_R0_clk;
  wire [7:0] mem_75_2_R0_data;
  wire  mem_75_2_R0_en;
  wire [25:0] mem_75_2_W0_addr;
  wire  mem_75_2_W0_clk;
  wire [7:0] mem_75_2_W0_data;
  wire  mem_75_2_W0_en;
  wire  mem_75_2_W0_mask;
  wire [25:0] mem_75_3_R0_addr;
  wire  mem_75_3_R0_clk;
  wire [7:0] mem_75_3_R0_data;
  wire  mem_75_3_R0_en;
  wire [25:0] mem_75_3_W0_addr;
  wire  mem_75_3_W0_clk;
  wire [7:0] mem_75_3_W0_data;
  wire  mem_75_3_W0_en;
  wire  mem_75_3_W0_mask;
  wire [25:0] mem_75_4_R0_addr;
  wire  mem_75_4_R0_clk;
  wire [7:0] mem_75_4_R0_data;
  wire  mem_75_4_R0_en;
  wire [25:0] mem_75_4_W0_addr;
  wire  mem_75_4_W0_clk;
  wire [7:0] mem_75_4_W0_data;
  wire  mem_75_4_W0_en;
  wire  mem_75_4_W0_mask;
  wire [25:0] mem_75_5_R0_addr;
  wire  mem_75_5_R0_clk;
  wire [7:0] mem_75_5_R0_data;
  wire  mem_75_5_R0_en;
  wire [25:0] mem_75_5_W0_addr;
  wire  mem_75_5_W0_clk;
  wire [7:0] mem_75_5_W0_data;
  wire  mem_75_5_W0_en;
  wire  mem_75_5_W0_mask;
  wire [25:0] mem_75_6_R0_addr;
  wire  mem_75_6_R0_clk;
  wire [7:0] mem_75_6_R0_data;
  wire  mem_75_6_R0_en;
  wire [25:0] mem_75_6_W0_addr;
  wire  mem_75_6_W0_clk;
  wire [7:0] mem_75_6_W0_data;
  wire  mem_75_6_W0_en;
  wire  mem_75_6_W0_mask;
  wire [25:0] mem_75_7_R0_addr;
  wire  mem_75_7_R0_clk;
  wire [7:0] mem_75_7_R0_data;
  wire  mem_75_7_R0_en;
  wire [25:0] mem_75_7_W0_addr;
  wire  mem_75_7_W0_clk;
  wire [7:0] mem_75_7_W0_data;
  wire  mem_75_7_W0_en;
  wire  mem_75_7_W0_mask;
  wire [25:0] mem_76_0_R0_addr;
  wire  mem_76_0_R0_clk;
  wire [7:0] mem_76_0_R0_data;
  wire  mem_76_0_R0_en;
  wire [25:0] mem_76_0_W0_addr;
  wire  mem_76_0_W0_clk;
  wire [7:0] mem_76_0_W0_data;
  wire  mem_76_0_W0_en;
  wire  mem_76_0_W0_mask;
  wire [25:0] mem_76_1_R0_addr;
  wire  mem_76_1_R0_clk;
  wire [7:0] mem_76_1_R0_data;
  wire  mem_76_1_R0_en;
  wire [25:0] mem_76_1_W0_addr;
  wire  mem_76_1_W0_clk;
  wire [7:0] mem_76_1_W0_data;
  wire  mem_76_1_W0_en;
  wire  mem_76_1_W0_mask;
  wire [25:0] mem_76_2_R0_addr;
  wire  mem_76_2_R0_clk;
  wire [7:0] mem_76_2_R0_data;
  wire  mem_76_2_R0_en;
  wire [25:0] mem_76_2_W0_addr;
  wire  mem_76_2_W0_clk;
  wire [7:0] mem_76_2_W0_data;
  wire  mem_76_2_W0_en;
  wire  mem_76_2_W0_mask;
  wire [25:0] mem_76_3_R0_addr;
  wire  mem_76_3_R0_clk;
  wire [7:0] mem_76_3_R0_data;
  wire  mem_76_3_R0_en;
  wire [25:0] mem_76_3_W0_addr;
  wire  mem_76_3_W0_clk;
  wire [7:0] mem_76_3_W0_data;
  wire  mem_76_3_W0_en;
  wire  mem_76_3_W0_mask;
  wire [25:0] mem_76_4_R0_addr;
  wire  mem_76_4_R0_clk;
  wire [7:0] mem_76_4_R0_data;
  wire  mem_76_4_R0_en;
  wire [25:0] mem_76_4_W0_addr;
  wire  mem_76_4_W0_clk;
  wire [7:0] mem_76_4_W0_data;
  wire  mem_76_4_W0_en;
  wire  mem_76_4_W0_mask;
  wire [25:0] mem_76_5_R0_addr;
  wire  mem_76_5_R0_clk;
  wire [7:0] mem_76_5_R0_data;
  wire  mem_76_5_R0_en;
  wire [25:0] mem_76_5_W0_addr;
  wire  mem_76_5_W0_clk;
  wire [7:0] mem_76_5_W0_data;
  wire  mem_76_5_W0_en;
  wire  mem_76_5_W0_mask;
  wire [25:0] mem_76_6_R0_addr;
  wire  mem_76_6_R0_clk;
  wire [7:0] mem_76_6_R0_data;
  wire  mem_76_6_R0_en;
  wire [25:0] mem_76_6_W0_addr;
  wire  mem_76_6_W0_clk;
  wire [7:0] mem_76_6_W0_data;
  wire  mem_76_6_W0_en;
  wire  mem_76_6_W0_mask;
  wire [25:0] mem_76_7_R0_addr;
  wire  mem_76_7_R0_clk;
  wire [7:0] mem_76_7_R0_data;
  wire  mem_76_7_R0_en;
  wire [25:0] mem_76_7_W0_addr;
  wire  mem_76_7_W0_clk;
  wire [7:0] mem_76_7_W0_data;
  wire  mem_76_7_W0_en;
  wire  mem_76_7_W0_mask;
  wire [25:0] mem_77_0_R0_addr;
  wire  mem_77_0_R0_clk;
  wire [7:0] mem_77_0_R0_data;
  wire  mem_77_0_R0_en;
  wire [25:0] mem_77_0_W0_addr;
  wire  mem_77_0_W0_clk;
  wire [7:0] mem_77_0_W0_data;
  wire  mem_77_0_W0_en;
  wire  mem_77_0_W0_mask;
  wire [25:0] mem_77_1_R0_addr;
  wire  mem_77_1_R0_clk;
  wire [7:0] mem_77_1_R0_data;
  wire  mem_77_1_R0_en;
  wire [25:0] mem_77_1_W0_addr;
  wire  mem_77_1_W0_clk;
  wire [7:0] mem_77_1_W0_data;
  wire  mem_77_1_W0_en;
  wire  mem_77_1_W0_mask;
  wire [25:0] mem_77_2_R0_addr;
  wire  mem_77_2_R0_clk;
  wire [7:0] mem_77_2_R0_data;
  wire  mem_77_2_R0_en;
  wire [25:0] mem_77_2_W0_addr;
  wire  mem_77_2_W0_clk;
  wire [7:0] mem_77_2_W0_data;
  wire  mem_77_2_W0_en;
  wire  mem_77_2_W0_mask;
  wire [25:0] mem_77_3_R0_addr;
  wire  mem_77_3_R0_clk;
  wire [7:0] mem_77_3_R0_data;
  wire  mem_77_3_R0_en;
  wire [25:0] mem_77_3_W0_addr;
  wire  mem_77_3_W0_clk;
  wire [7:0] mem_77_3_W0_data;
  wire  mem_77_3_W0_en;
  wire  mem_77_3_W0_mask;
  wire [25:0] mem_77_4_R0_addr;
  wire  mem_77_4_R0_clk;
  wire [7:0] mem_77_4_R0_data;
  wire  mem_77_4_R0_en;
  wire [25:0] mem_77_4_W0_addr;
  wire  mem_77_4_W0_clk;
  wire [7:0] mem_77_4_W0_data;
  wire  mem_77_4_W0_en;
  wire  mem_77_4_W0_mask;
  wire [25:0] mem_77_5_R0_addr;
  wire  mem_77_5_R0_clk;
  wire [7:0] mem_77_5_R0_data;
  wire  mem_77_5_R0_en;
  wire [25:0] mem_77_5_W0_addr;
  wire  mem_77_5_W0_clk;
  wire [7:0] mem_77_5_W0_data;
  wire  mem_77_5_W0_en;
  wire  mem_77_5_W0_mask;
  wire [25:0] mem_77_6_R0_addr;
  wire  mem_77_6_R0_clk;
  wire [7:0] mem_77_6_R0_data;
  wire  mem_77_6_R0_en;
  wire [25:0] mem_77_6_W0_addr;
  wire  mem_77_6_W0_clk;
  wire [7:0] mem_77_6_W0_data;
  wire  mem_77_6_W0_en;
  wire  mem_77_6_W0_mask;
  wire [25:0] mem_77_7_R0_addr;
  wire  mem_77_7_R0_clk;
  wire [7:0] mem_77_7_R0_data;
  wire  mem_77_7_R0_en;
  wire [25:0] mem_77_7_W0_addr;
  wire  mem_77_7_W0_clk;
  wire [7:0] mem_77_7_W0_data;
  wire  mem_77_7_W0_en;
  wire  mem_77_7_W0_mask;
  wire [25:0] mem_78_0_R0_addr;
  wire  mem_78_0_R0_clk;
  wire [7:0] mem_78_0_R0_data;
  wire  mem_78_0_R0_en;
  wire [25:0] mem_78_0_W0_addr;
  wire  mem_78_0_W0_clk;
  wire [7:0] mem_78_0_W0_data;
  wire  mem_78_0_W0_en;
  wire  mem_78_0_W0_mask;
  wire [25:0] mem_78_1_R0_addr;
  wire  mem_78_1_R0_clk;
  wire [7:0] mem_78_1_R0_data;
  wire  mem_78_1_R0_en;
  wire [25:0] mem_78_1_W0_addr;
  wire  mem_78_1_W0_clk;
  wire [7:0] mem_78_1_W0_data;
  wire  mem_78_1_W0_en;
  wire  mem_78_1_W0_mask;
  wire [25:0] mem_78_2_R0_addr;
  wire  mem_78_2_R0_clk;
  wire [7:0] mem_78_2_R0_data;
  wire  mem_78_2_R0_en;
  wire [25:0] mem_78_2_W0_addr;
  wire  mem_78_2_W0_clk;
  wire [7:0] mem_78_2_W0_data;
  wire  mem_78_2_W0_en;
  wire  mem_78_2_W0_mask;
  wire [25:0] mem_78_3_R0_addr;
  wire  mem_78_3_R0_clk;
  wire [7:0] mem_78_3_R0_data;
  wire  mem_78_3_R0_en;
  wire [25:0] mem_78_3_W0_addr;
  wire  mem_78_3_W0_clk;
  wire [7:0] mem_78_3_W0_data;
  wire  mem_78_3_W0_en;
  wire  mem_78_3_W0_mask;
  wire [25:0] mem_78_4_R0_addr;
  wire  mem_78_4_R0_clk;
  wire [7:0] mem_78_4_R0_data;
  wire  mem_78_4_R0_en;
  wire [25:0] mem_78_4_W0_addr;
  wire  mem_78_4_W0_clk;
  wire [7:0] mem_78_4_W0_data;
  wire  mem_78_4_W0_en;
  wire  mem_78_4_W0_mask;
  wire [25:0] mem_78_5_R0_addr;
  wire  mem_78_5_R0_clk;
  wire [7:0] mem_78_5_R0_data;
  wire  mem_78_5_R0_en;
  wire [25:0] mem_78_5_W0_addr;
  wire  mem_78_5_W0_clk;
  wire [7:0] mem_78_5_W0_data;
  wire  mem_78_5_W0_en;
  wire  mem_78_5_W0_mask;
  wire [25:0] mem_78_6_R0_addr;
  wire  mem_78_6_R0_clk;
  wire [7:0] mem_78_6_R0_data;
  wire  mem_78_6_R0_en;
  wire [25:0] mem_78_6_W0_addr;
  wire  mem_78_6_W0_clk;
  wire [7:0] mem_78_6_W0_data;
  wire  mem_78_6_W0_en;
  wire  mem_78_6_W0_mask;
  wire [25:0] mem_78_7_R0_addr;
  wire  mem_78_7_R0_clk;
  wire [7:0] mem_78_7_R0_data;
  wire  mem_78_7_R0_en;
  wire [25:0] mem_78_7_W0_addr;
  wire  mem_78_7_W0_clk;
  wire [7:0] mem_78_7_W0_data;
  wire  mem_78_7_W0_en;
  wire  mem_78_7_W0_mask;
  wire [25:0] mem_79_0_R0_addr;
  wire  mem_79_0_R0_clk;
  wire [7:0] mem_79_0_R0_data;
  wire  mem_79_0_R0_en;
  wire [25:0] mem_79_0_W0_addr;
  wire  mem_79_0_W0_clk;
  wire [7:0] mem_79_0_W0_data;
  wire  mem_79_0_W0_en;
  wire  mem_79_0_W0_mask;
  wire [25:0] mem_79_1_R0_addr;
  wire  mem_79_1_R0_clk;
  wire [7:0] mem_79_1_R0_data;
  wire  mem_79_1_R0_en;
  wire [25:0] mem_79_1_W0_addr;
  wire  mem_79_1_W0_clk;
  wire [7:0] mem_79_1_W0_data;
  wire  mem_79_1_W0_en;
  wire  mem_79_1_W0_mask;
  wire [25:0] mem_79_2_R0_addr;
  wire  mem_79_2_R0_clk;
  wire [7:0] mem_79_2_R0_data;
  wire  mem_79_2_R0_en;
  wire [25:0] mem_79_2_W0_addr;
  wire  mem_79_2_W0_clk;
  wire [7:0] mem_79_2_W0_data;
  wire  mem_79_2_W0_en;
  wire  mem_79_2_W0_mask;
  wire [25:0] mem_79_3_R0_addr;
  wire  mem_79_3_R0_clk;
  wire [7:0] mem_79_3_R0_data;
  wire  mem_79_3_R0_en;
  wire [25:0] mem_79_3_W0_addr;
  wire  mem_79_3_W0_clk;
  wire [7:0] mem_79_3_W0_data;
  wire  mem_79_3_W0_en;
  wire  mem_79_3_W0_mask;
  wire [25:0] mem_79_4_R0_addr;
  wire  mem_79_4_R0_clk;
  wire [7:0] mem_79_4_R0_data;
  wire  mem_79_4_R0_en;
  wire [25:0] mem_79_4_W0_addr;
  wire  mem_79_4_W0_clk;
  wire [7:0] mem_79_4_W0_data;
  wire  mem_79_4_W0_en;
  wire  mem_79_4_W0_mask;
  wire [25:0] mem_79_5_R0_addr;
  wire  mem_79_5_R0_clk;
  wire [7:0] mem_79_5_R0_data;
  wire  mem_79_5_R0_en;
  wire [25:0] mem_79_5_W0_addr;
  wire  mem_79_5_W0_clk;
  wire [7:0] mem_79_5_W0_data;
  wire  mem_79_5_W0_en;
  wire  mem_79_5_W0_mask;
  wire [25:0] mem_79_6_R0_addr;
  wire  mem_79_6_R0_clk;
  wire [7:0] mem_79_6_R0_data;
  wire  mem_79_6_R0_en;
  wire [25:0] mem_79_6_W0_addr;
  wire  mem_79_6_W0_clk;
  wire [7:0] mem_79_6_W0_data;
  wire  mem_79_6_W0_en;
  wire  mem_79_6_W0_mask;
  wire [25:0] mem_79_7_R0_addr;
  wire  mem_79_7_R0_clk;
  wire [7:0] mem_79_7_R0_data;
  wire  mem_79_7_R0_en;
  wire [25:0] mem_79_7_W0_addr;
  wire  mem_79_7_W0_clk;
  wire [7:0] mem_79_7_W0_data;
  wire  mem_79_7_W0_en;
  wire  mem_79_7_W0_mask;
  wire [25:0] mem_80_0_R0_addr;
  wire  mem_80_0_R0_clk;
  wire [7:0] mem_80_0_R0_data;
  wire  mem_80_0_R0_en;
  wire [25:0] mem_80_0_W0_addr;
  wire  mem_80_0_W0_clk;
  wire [7:0] mem_80_0_W0_data;
  wire  mem_80_0_W0_en;
  wire  mem_80_0_W0_mask;
  wire [25:0] mem_80_1_R0_addr;
  wire  mem_80_1_R0_clk;
  wire [7:0] mem_80_1_R0_data;
  wire  mem_80_1_R0_en;
  wire [25:0] mem_80_1_W0_addr;
  wire  mem_80_1_W0_clk;
  wire [7:0] mem_80_1_W0_data;
  wire  mem_80_1_W0_en;
  wire  mem_80_1_W0_mask;
  wire [25:0] mem_80_2_R0_addr;
  wire  mem_80_2_R0_clk;
  wire [7:0] mem_80_2_R0_data;
  wire  mem_80_2_R0_en;
  wire [25:0] mem_80_2_W0_addr;
  wire  mem_80_2_W0_clk;
  wire [7:0] mem_80_2_W0_data;
  wire  mem_80_2_W0_en;
  wire  mem_80_2_W0_mask;
  wire [25:0] mem_80_3_R0_addr;
  wire  mem_80_3_R0_clk;
  wire [7:0] mem_80_3_R0_data;
  wire  mem_80_3_R0_en;
  wire [25:0] mem_80_3_W0_addr;
  wire  mem_80_3_W0_clk;
  wire [7:0] mem_80_3_W0_data;
  wire  mem_80_3_W0_en;
  wire  mem_80_3_W0_mask;
  wire [25:0] mem_80_4_R0_addr;
  wire  mem_80_4_R0_clk;
  wire [7:0] mem_80_4_R0_data;
  wire  mem_80_4_R0_en;
  wire [25:0] mem_80_4_W0_addr;
  wire  mem_80_4_W0_clk;
  wire [7:0] mem_80_4_W0_data;
  wire  mem_80_4_W0_en;
  wire  mem_80_4_W0_mask;
  wire [25:0] mem_80_5_R0_addr;
  wire  mem_80_5_R0_clk;
  wire [7:0] mem_80_5_R0_data;
  wire  mem_80_5_R0_en;
  wire [25:0] mem_80_5_W0_addr;
  wire  mem_80_5_W0_clk;
  wire [7:0] mem_80_5_W0_data;
  wire  mem_80_5_W0_en;
  wire  mem_80_5_W0_mask;
  wire [25:0] mem_80_6_R0_addr;
  wire  mem_80_6_R0_clk;
  wire [7:0] mem_80_6_R0_data;
  wire  mem_80_6_R0_en;
  wire [25:0] mem_80_6_W0_addr;
  wire  mem_80_6_W0_clk;
  wire [7:0] mem_80_6_W0_data;
  wire  mem_80_6_W0_en;
  wire  mem_80_6_W0_mask;
  wire [25:0] mem_80_7_R0_addr;
  wire  mem_80_7_R0_clk;
  wire [7:0] mem_80_7_R0_data;
  wire  mem_80_7_R0_en;
  wire [25:0] mem_80_7_W0_addr;
  wire  mem_80_7_W0_clk;
  wire [7:0] mem_80_7_W0_data;
  wire  mem_80_7_W0_en;
  wire  mem_80_7_W0_mask;
  wire [25:0] mem_81_0_R0_addr;
  wire  mem_81_0_R0_clk;
  wire [7:0] mem_81_0_R0_data;
  wire  mem_81_0_R0_en;
  wire [25:0] mem_81_0_W0_addr;
  wire  mem_81_0_W0_clk;
  wire [7:0] mem_81_0_W0_data;
  wire  mem_81_0_W0_en;
  wire  mem_81_0_W0_mask;
  wire [25:0] mem_81_1_R0_addr;
  wire  mem_81_1_R0_clk;
  wire [7:0] mem_81_1_R0_data;
  wire  mem_81_1_R0_en;
  wire [25:0] mem_81_1_W0_addr;
  wire  mem_81_1_W0_clk;
  wire [7:0] mem_81_1_W0_data;
  wire  mem_81_1_W0_en;
  wire  mem_81_1_W0_mask;
  wire [25:0] mem_81_2_R0_addr;
  wire  mem_81_2_R0_clk;
  wire [7:0] mem_81_2_R0_data;
  wire  mem_81_2_R0_en;
  wire [25:0] mem_81_2_W0_addr;
  wire  mem_81_2_W0_clk;
  wire [7:0] mem_81_2_W0_data;
  wire  mem_81_2_W0_en;
  wire  mem_81_2_W0_mask;
  wire [25:0] mem_81_3_R0_addr;
  wire  mem_81_3_R0_clk;
  wire [7:0] mem_81_3_R0_data;
  wire  mem_81_3_R0_en;
  wire [25:0] mem_81_3_W0_addr;
  wire  mem_81_3_W0_clk;
  wire [7:0] mem_81_3_W0_data;
  wire  mem_81_3_W0_en;
  wire  mem_81_3_W0_mask;
  wire [25:0] mem_81_4_R0_addr;
  wire  mem_81_4_R0_clk;
  wire [7:0] mem_81_4_R0_data;
  wire  mem_81_4_R0_en;
  wire [25:0] mem_81_4_W0_addr;
  wire  mem_81_4_W0_clk;
  wire [7:0] mem_81_4_W0_data;
  wire  mem_81_4_W0_en;
  wire  mem_81_4_W0_mask;
  wire [25:0] mem_81_5_R0_addr;
  wire  mem_81_5_R0_clk;
  wire [7:0] mem_81_5_R0_data;
  wire  mem_81_5_R0_en;
  wire [25:0] mem_81_5_W0_addr;
  wire  mem_81_5_W0_clk;
  wire [7:0] mem_81_5_W0_data;
  wire  mem_81_5_W0_en;
  wire  mem_81_5_W0_mask;
  wire [25:0] mem_81_6_R0_addr;
  wire  mem_81_6_R0_clk;
  wire [7:0] mem_81_6_R0_data;
  wire  mem_81_6_R0_en;
  wire [25:0] mem_81_6_W0_addr;
  wire  mem_81_6_W0_clk;
  wire [7:0] mem_81_6_W0_data;
  wire  mem_81_6_W0_en;
  wire  mem_81_6_W0_mask;
  wire [25:0] mem_81_7_R0_addr;
  wire  mem_81_7_R0_clk;
  wire [7:0] mem_81_7_R0_data;
  wire  mem_81_7_R0_en;
  wire [25:0] mem_81_7_W0_addr;
  wire  mem_81_7_W0_clk;
  wire [7:0] mem_81_7_W0_data;
  wire  mem_81_7_W0_en;
  wire  mem_81_7_W0_mask;
  wire [25:0] mem_82_0_R0_addr;
  wire  mem_82_0_R0_clk;
  wire [7:0] mem_82_0_R0_data;
  wire  mem_82_0_R0_en;
  wire [25:0] mem_82_0_W0_addr;
  wire  mem_82_0_W0_clk;
  wire [7:0] mem_82_0_W0_data;
  wire  mem_82_0_W0_en;
  wire  mem_82_0_W0_mask;
  wire [25:0] mem_82_1_R0_addr;
  wire  mem_82_1_R0_clk;
  wire [7:0] mem_82_1_R0_data;
  wire  mem_82_1_R0_en;
  wire [25:0] mem_82_1_W0_addr;
  wire  mem_82_1_W0_clk;
  wire [7:0] mem_82_1_W0_data;
  wire  mem_82_1_W0_en;
  wire  mem_82_1_W0_mask;
  wire [25:0] mem_82_2_R0_addr;
  wire  mem_82_2_R0_clk;
  wire [7:0] mem_82_2_R0_data;
  wire  mem_82_2_R0_en;
  wire [25:0] mem_82_2_W0_addr;
  wire  mem_82_2_W0_clk;
  wire [7:0] mem_82_2_W0_data;
  wire  mem_82_2_W0_en;
  wire  mem_82_2_W0_mask;
  wire [25:0] mem_82_3_R0_addr;
  wire  mem_82_3_R0_clk;
  wire [7:0] mem_82_3_R0_data;
  wire  mem_82_3_R0_en;
  wire [25:0] mem_82_3_W0_addr;
  wire  mem_82_3_W0_clk;
  wire [7:0] mem_82_3_W0_data;
  wire  mem_82_3_W0_en;
  wire  mem_82_3_W0_mask;
  wire [25:0] mem_82_4_R0_addr;
  wire  mem_82_4_R0_clk;
  wire [7:0] mem_82_4_R0_data;
  wire  mem_82_4_R0_en;
  wire [25:0] mem_82_4_W0_addr;
  wire  mem_82_4_W0_clk;
  wire [7:0] mem_82_4_W0_data;
  wire  mem_82_4_W0_en;
  wire  mem_82_4_W0_mask;
  wire [25:0] mem_82_5_R0_addr;
  wire  mem_82_5_R0_clk;
  wire [7:0] mem_82_5_R0_data;
  wire  mem_82_5_R0_en;
  wire [25:0] mem_82_5_W0_addr;
  wire  mem_82_5_W0_clk;
  wire [7:0] mem_82_5_W0_data;
  wire  mem_82_5_W0_en;
  wire  mem_82_5_W0_mask;
  wire [25:0] mem_82_6_R0_addr;
  wire  mem_82_6_R0_clk;
  wire [7:0] mem_82_6_R0_data;
  wire  mem_82_6_R0_en;
  wire [25:0] mem_82_6_W0_addr;
  wire  mem_82_6_W0_clk;
  wire [7:0] mem_82_6_W0_data;
  wire  mem_82_6_W0_en;
  wire  mem_82_6_W0_mask;
  wire [25:0] mem_82_7_R0_addr;
  wire  mem_82_7_R0_clk;
  wire [7:0] mem_82_7_R0_data;
  wire  mem_82_7_R0_en;
  wire [25:0] mem_82_7_W0_addr;
  wire  mem_82_7_W0_clk;
  wire [7:0] mem_82_7_W0_data;
  wire  mem_82_7_W0_en;
  wire  mem_82_7_W0_mask;
  wire [25:0] mem_83_0_R0_addr;
  wire  mem_83_0_R0_clk;
  wire [7:0] mem_83_0_R0_data;
  wire  mem_83_0_R0_en;
  wire [25:0] mem_83_0_W0_addr;
  wire  mem_83_0_W0_clk;
  wire [7:0] mem_83_0_W0_data;
  wire  mem_83_0_W0_en;
  wire  mem_83_0_W0_mask;
  wire [25:0] mem_83_1_R0_addr;
  wire  mem_83_1_R0_clk;
  wire [7:0] mem_83_1_R0_data;
  wire  mem_83_1_R0_en;
  wire [25:0] mem_83_1_W0_addr;
  wire  mem_83_1_W0_clk;
  wire [7:0] mem_83_1_W0_data;
  wire  mem_83_1_W0_en;
  wire  mem_83_1_W0_mask;
  wire [25:0] mem_83_2_R0_addr;
  wire  mem_83_2_R0_clk;
  wire [7:0] mem_83_2_R0_data;
  wire  mem_83_2_R0_en;
  wire [25:0] mem_83_2_W0_addr;
  wire  mem_83_2_W0_clk;
  wire [7:0] mem_83_2_W0_data;
  wire  mem_83_2_W0_en;
  wire  mem_83_2_W0_mask;
  wire [25:0] mem_83_3_R0_addr;
  wire  mem_83_3_R0_clk;
  wire [7:0] mem_83_3_R0_data;
  wire  mem_83_3_R0_en;
  wire [25:0] mem_83_3_W0_addr;
  wire  mem_83_3_W0_clk;
  wire [7:0] mem_83_3_W0_data;
  wire  mem_83_3_W0_en;
  wire  mem_83_3_W0_mask;
  wire [25:0] mem_83_4_R0_addr;
  wire  mem_83_4_R0_clk;
  wire [7:0] mem_83_4_R0_data;
  wire  mem_83_4_R0_en;
  wire [25:0] mem_83_4_W0_addr;
  wire  mem_83_4_W0_clk;
  wire [7:0] mem_83_4_W0_data;
  wire  mem_83_4_W0_en;
  wire  mem_83_4_W0_mask;
  wire [25:0] mem_83_5_R0_addr;
  wire  mem_83_5_R0_clk;
  wire [7:0] mem_83_5_R0_data;
  wire  mem_83_5_R0_en;
  wire [25:0] mem_83_5_W0_addr;
  wire  mem_83_5_W0_clk;
  wire [7:0] mem_83_5_W0_data;
  wire  mem_83_5_W0_en;
  wire  mem_83_5_W0_mask;
  wire [25:0] mem_83_6_R0_addr;
  wire  mem_83_6_R0_clk;
  wire [7:0] mem_83_6_R0_data;
  wire  mem_83_6_R0_en;
  wire [25:0] mem_83_6_W0_addr;
  wire  mem_83_6_W0_clk;
  wire [7:0] mem_83_6_W0_data;
  wire  mem_83_6_W0_en;
  wire  mem_83_6_W0_mask;
  wire [25:0] mem_83_7_R0_addr;
  wire  mem_83_7_R0_clk;
  wire [7:0] mem_83_7_R0_data;
  wire  mem_83_7_R0_en;
  wire [25:0] mem_83_7_W0_addr;
  wire  mem_83_7_W0_clk;
  wire [7:0] mem_83_7_W0_data;
  wire  mem_83_7_W0_en;
  wire  mem_83_7_W0_mask;
  wire [25:0] mem_84_0_R0_addr;
  wire  mem_84_0_R0_clk;
  wire [7:0] mem_84_0_R0_data;
  wire  mem_84_0_R0_en;
  wire [25:0] mem_84_0_W0_addr;
  wire  mem_84_0_W0_clk;
  wire [7:0] mem_84_0_W0_data;
  wire  mem_84_0_W0_en;
  wire  mem_84_0_W0_mask;
  wire [25:0] mem_84_1_R0_addr;
  wire  mem_84_1_R0_clk;
  wire [7:0] mem_84_1_R0_data;
  wire  mem_84_1_R0_en;
  wire [25:0] mem_84_1_W0_addr;
  wire  mem_84_1_W0_clk;
  wire [7:0] mem_84_1_W0_data;
  wire  mem_84_1_W0_en;
  wire  mem_84_1_W0_mask;
  wire [25:0] mem_84_2_R0_addr;
  wire  mem_84_2_R0_clk;
  wire [7:0] mem_84_2_R0_data;
  wire  mem_84_2_R0_en;
  wire [25:0] mem_84_2_W0_addr;
  wire  mem_84_2_W0_clk;
  wire [7:0] mem_84_2_W0_data;
  wire  mem_84_2_W0_en;
  wire  mem_84_2_W0_mask;
  wire [25:0] mem_84_3_R0_addr;
  wire  mem_84_3_R0_clk;
  wire [7:0] mem_84_3_R0_data;
  wire  mem_84_3_R0_en;
  wire [25:0] mem_84_3_W0_addr;
  wire  mem_84_3_W0_clk;
  wire [7:0] mem_84_3_W0_data;
  wire  mem_84_3_W0_en;
  wire  mem_84_3_W0_mask;
  wire [25:0] mem_84_4_R0_addr;
  wire  mem_84_4_R0_clk;
  wire [7:0] mem_84_4_R0_data;
  wire  mem_84_4_R0_en;
  wire [25:0] mem_84_4_W0_addr;
  wire  mem_84_4_W0_clk;
  wire [7:0] mem_84_4_W0_data;
  wire  mem_84_4_W0_en;
  wire  mem_84_4_W0_mask;
  wire [25:0] mem_84_5_R0_addr;
  wire  mem_84_5_R0_clk;
  wire [7:0] mem_84_5_R0_data;
  wire  mem_84_5_R0_en;
  wire [25:0] mem_84_5_W0_addr;
  wire  mem_84_5_W0_clk;
  wire [7:0] mem_84_5_W0_data;
  wire  mem_84_5_W0_en;
  wire  mem_84_5_W0_mask;
  wire [25:0] mem_84_6_R0_addr;
  wire  mem_84_6_R0_clk;
  wire [7:0] mem_84_6_R0_data;
  wire  mem_84_6_R0_en;
  wire [25:0] mem_84_6_W0_addr;
  wire  mem_84_6_W0_clk;
  wire [7:0] mem_84_6_W0_data;
  wire  mem_84_6_W0_en;
  wire  mem_84_6_W0_mask;
  wire [25:0] mem_84_7_R0_addr;
  wire  mem_84_7_R0_clk;
  wire [7:0] mem_84_7_R0_data;
  wire  mem_84_7_R0_en;
  wire [25:0] mem_84_7_W0_addr;
  wire  mem_84_7_W0_clk;
  wire [7:0] mem_84_7_W0_data;
  wire  mem_84_7_W0_en;
  wire  mem_84_7_W0_mask;
  wire [25:0] mem_85_0_R0_addr;
  wire  mem_85_0_R0_clk;
  wire [7:0] mem_85_0_R0_data;
  wire  mem_85_0_R0_en;
  wire [25:0] mem_85_0_W0_addr;
  wire  mem_85_0_W0_clk;
  wire [7:0] mem_85_0_W0_data;
  wire  mem_85_0_W0_en;
  wire  mem_85_0_W0_mask;
  wire [25:0] mem_85_1_R0_addr;
  wire  mem_85_1_R0_clk;
  wire [7:0] mem_85_1_R0_data;
  wire  mem_85_1_R0_en;
  wire [25:0] mem_85_1_W0_addr;
  wire  mem_85_1_W0_clk;
  wire [7:0] mem_85_1_W0_data;
  wire  mem_85_1_W0_en;
  wire  mem_85_1_W0_mask;
  wire [25:0] mem_85_2_R0_addr;
  wire  mem_85_2_R0_clk;
  wire [7:0] mem_85_2_R0_data;
  wire  mem_85_2_R0_en;
  wire [25:0] mem_85_2_W0_addr;
  wire  mem_85_2_W0_clk;
  wire [7:0] mem_85_2_W0_data;
  wire  mem_85_2_W0_en;
  wire  mem_85_2_W0_mask;
  wire [25:0] mem_85_3_R0_addr;
  wire  mem_85_3_R0_clk;
  wire [7:0] mem_85_3_R0_data;
  wire  mem_85_3_R0_en;
  wire [25:0] mem_85_3_W0_addr;
  wire  mem_85_3_W0_clk;
  wire [7:0] mem_85_3_W0_data;
  wire  mem_85_3_W0_en;
  wire  mem_85_3_W0_mask;
  wire [25:0] mem_85_4_R0_addr;
  wire  mem_85_4_R0_clk;
  wire [7:0] mem_85_4_R0_data;
  wire  mem_85_4_R0_en;
  wire [25:0] mem_85_4_W0_addr;
  wire  mem_85_4_W0_clk;
  wire [7:0] mem_85_4_W0_data;
  wire  mem_85_4_W0_en;
  wire  mem_85_4_W0_mask;
  wire [25:0] mem_85_5_R0_addr;
  wire  mem_85_5_R0_clk;
  wire [7:0] mem_85_5_R0_data;
  wire  mem_85_5_R0_en;
  wire [25:0] mem_85_5_W0_addr;
  wire  mem_85_5_W0_clk;
  wire [7:0] mem_85_5_W0_data;
  wire  mem_85_5_W0_en;
  wire  mem_85_5_W0_mask;
  wire [25:0] mem_85_6_R0_addr;
  wire  mem_85_6_R0_clk;
  wire [7:0] mem_85_6_R0_data;
  wire  mem_85_6_R0_en;
  wire [25:0] mem_85_6_W0_addr;
  wire  mem_85_6_W0_clk;
  wire [7:0] mem_85_6_W0_data;
  wire  mem_85_6_W0_en;
  wire  mem_85_6_W0_mask;
  wire [25:0] mem_85_7_R0_addr;
  wire  mem_85_7_R0_clk;
  wire [7:0] mem_85_7_R0_data;
  wire  mem_85_7_R0_en;
  wire [25:0] mem_85_7_W0_addr;
  wire  mem_85_7_W0_clk;
  wire [7:0] mem_85_7_W0_data;
  wire  mem_85_7_W0_en;
  wire  mem_85_7_W0_mask;
  wire [25:0] mem_86_0_R0_addr;
  wire  mem_86_0_R0_clk;
  wire [7:0] mem_86_0_R0_data;
  wire  mem_86_0_R0_en;
  wire [25:0] mem_86_0_W0_addr;
  wire  mem_86_0_W0_clk;
  wire [7:0] mem_86_0_W0_data;
  wire  mem_86_0_W0_en;
  wire  mem_86_0_W0_mask;
  wire [25:0] mem_86_1_R0_addr;
  wire  mem_86_1_R0_clk;
  wire [7:0] mem_86_1_R0_data;
  wire  mem_86_1_R0_en;
  wire [25:0] mem_86_1_W0_addr;
  wire  mem_86_1_W0_clk;
  wire [7:0] mem_86_1_W0_data;
  wire  mem_86_1_W0_en;
  wire  mem_86_1_W0_mask;
  wire [25:0] mem_86_2_R0_addr;
  wire  mem_86_2_R0_clk;
  wire [7:0] mem_86_2_R0_data;
  wire  mem_86_2_R0_en;
  wire [25:0] mem_86_2_W0_addr;
  wire  mem_86_2_W0_clk;
  wire [7:0] mem_86_2_W0_data;
  wire  mem_86_2_W0_en;
  wire  mem_86_2_W0_mask;
  wire [25:0] mem_86_3_R0_addr;
  wire  mem_86_3_R0_clk;
  wire [7:0] mem_86_3_R0_data;
  wire  mem_86_3_R0_en;
  wire [25:0] mem_86_3_W0_addr;
  wire  mem_86_3_W0_clk;
  wire [7:0] mem_86_3_W0_data;
  wire  mem_86_3_W0_en;
  wire  mem_86_3_W0_mask;
  wire [25:0] mem_86_4_R0_addr;
  wire  mem_86_4_R0_clk;
  wire [7:0] mem_86_4_R0_data;
  wire  mem_86_4_R0_en;
  wire [25:0] mem_86_4_W0_addr;
  wire  mem_86_4_W0_clk;
  wire [7:0] mem_86_4_W0_data;
  wire  mem_86_4_W0_en;
  wire  mem_86_4_W0_mask;
  wire [25:0] mem_86_5_R0_addr;
  wire  mem_86_5_R0_clk;
  wire [7:0] mem_86_5_R0_data;
  wire  mem_86_5_R0_en;
  wire [25:0] mem_86_5_W0_addr;
  wire  mem_86_5_W0_clk;
  wire [7:0] mem_86_5_W0_data;
  wire  mem_86_5_W0_en;
  wire  mem_86_5_W0_mask;
  wire [25:0] mem_86_6_R0_addr;
  wire  mem_86_6_R0_clk;
  wire [7:0] mem_86_6_R0_data;
  wire  mem_86_6_R0_en;
  wire [25:0] mem_86_6_W0_addr;
  wire  mem_86_6_W0_clk;
  wire [7:0] mem_86_6_W0_data;
  wire  mem_86_6_W0_en;
  wire  mem_86_6_W0_mask;
  wire [25:0] mem_86_7_R0_addr;
  wire  mem_86_7_R0_clk;
  wire [7:0] mem_86_7_R0_data;
  wire  mem_86_7_R0_en;
  wire [25:0] mem_86_7_W0_addr;
  wire  mem_86_7_W0_clk;
  wire [7:0] mem_86_7_W0_data;
  wire  mem_86_7_W0_en;
  wire  mem_86_7_W0_mask;
  wire [25:0] mem_87_0_R0_addr;
  wire  mem_87_0_R0_clk;
  wire [7:0] mem_87_0_R0_data;
  wire  mem_87_0_R0_en;
  wire [25:0] mem_87_0_W0_addr;
  wire  mem_87_0_W0_clk;
  wire [7:0] mem_87_0_W0_data;
  wire  mem_87_0_W0_en;
  wire  mem_87_0_W0_mask;
  wire [25:0] mem_87_1_R0_addr;
  wire  mem_87_1_R0_clk;
  wire [7:0] mem_87_1_R0_data;
  wire  mem_87_1_R0_en;
  wire [25:0] mem_87_1_W0_addr;
  wire  mem_87_1_W0_clk;
  wire [7:0] mem_87_1_W0_data;
  wire  mem_87_1_W0_en;
  wire  mem_87_1_W0_mask;
  wire [25:0] mem_87_2_R0_addr;
  wire  mem_87_2_R0_clk;
  wire [7:0] mem_87_2_R0_data;
  wire  mem_87_2_R0_en;
  wire [25:0] mem_87_2_W0_addr;
  wire  mem_87_2_W0_clk;
  wire [7:0] mem_87_2_W0_data;
  wire  mem_87_2_W0_en;
  wire  mem_87_2_W0_mask;
  wire [25:0] mem_87_3_R0_addr;
  wire  mem_87_3_R0_clk;
  wire [7:0] mem_87_3_R0_data;
  wire  mem_87_3_R0_en;
  wire [25:0] mem_87_3_W0_addr;
  wire  mem_87_3_W0_clk;
  wire [7:0] mem_87_3_W0_data;
  wire  mem_87_3_W0_en;
  wire  mem_87_3_W0_mask;
  wire [25:0] mem_87_4_R0_addr;
  wire  mem_87_4_R0_clk;
  wire [7:0] mem_87_4_R0_data;
  wire  mem_87_4_R0_en;
  wire [25:0] mem_87_4_W0_addr;
  wire  mem_87_4_W0_clk;
  wire [7:0] mem_87_4_W0_data;
  wire  mem_87_4_W0_en;
  wire  mem_87_4_W0_mask;
  wire [25:0] mem_87_5_R0_addr;
  wire  mem_87_5_R0_clk;
  wire [7:0] mem_87_5_R0_data;
  wire  mem_87_5_R0_en;
  wire [25:0] mem_87_5_W0_addr;
  wire  mem_87_5_W0_clk;
  wire [7:0] mem_87_5_W0_data;
  wire  mem_87_5_W0_en;
  wire  mem_87_5_W0_mask;
  wire [25:0] mem_87_6_R0_addr;
  wire  mem_87_6_R0_clk;
  wire [7:0] mem_87_6_R0_data;
  wire  mem_87_6_R0_en;
  wire [25:0] mem_87_6_W0_addr;
  wire  mem_87_6_W0_clk;
  wire [7:0] mem_87_6_W0_data;
  wire  mem_87_6_W0_en;
  wire  mem_87_6_W0_mask;
  wire [25:0] mem_87_7_R0_addr;
  wire  mem_87_7_R0_clk;
  wire [7:0] mem_87_7_R0_data;
  wire  mem_87_7_R0_en;
  wire [25:0] mem_87_7_W0_addr;
  wire  mem_87_7_W0_clk;
  wire [7:0] mem_87_7_W0_data;
  wire  mem_87_7_W0_en;
  wire  mem_87_7_W0_mask;
  wire [25:0] mem_88_0_R0_addr;
  wire  mem_88_0_R0_clk;
  wire [7:0] mem_88_0_R0_data;
  wire  mem_88_0_R0_en;
  wire [25:0] mem_88_0_W0_addr;
  wire  mem_88_0_W0_clk;
  wire [7:0] mem_88_0_W0_data;
  wire  mem_88_0_W0_en;
  wire  mem_88_0_W0_mask;
  wire [25:0] mem_88_1_R0_addr;
  wire  mem_88_1_R0_clk;
  wire [7:0] mem_88_1_R0_data;
  wire  mem_88_1_R0_en;
  wire [25:0] mem_88_1_W0_addr;
  wire  mem_88_1_W0_clk;
  wire [7:0] mem_88_1_W0_data;
  wire  mem_88_1_W0_en;
  wire  mem_88_1_W0_mask;
  wire [25:0] mem_88_2_R0_addr;
  wire  mem_88_2_R0_clk;
  wire [7:0] mem_88_2_R0_data;
  wire  mem_88_2_R0_en;
  wire [25:0] mem_88_2_W0_addr;
  wire  mem_88_2_W0_clk;
  wire [7:0] mem_88_2_W0_data;
  wire  mem_88_2_W0_en;
  wire  mem_88_2_W0_mask;
  wire [25:0] mem_88_3_R0_addr;
  wire  mem_88_3_R0_clk;
  wire [7:0] mem_88_3_R0_data;
  wire  mem_88_3_R0_en;
  wire [25:0] mem_88_3_W0_addr;
  wire  mem_88_3_W0_clk;
  wire [7:0] mem_88_3_W0_data;
  wire  mem_88_3_W0_en;
  wire  mem_88_3_W0_mask;
  wire [25:0] mem_88_4_R0_addr;
  wire  mem_88_4_R0_clk;
  wire [7:0] mem_88_4_R0_data;
  wire  mem_88_4_R0_en;
  wire [25:0] mem_88_4_W0_addr;
  wire  mem_88_4_W0_clk;
  wire [7:0] mem_88_4_W0_data;
  wire  mem_88_4_W0_en;
  wire  mem_88_4_W0_mask;
  wire [25:0] mem_88_5_R0_addr;
  wire  mem_88_5_R0_clk;
  wire [7:0] mem_88_5_R0_data;
  wire  mem_88_5_R0_en;
  wire [25:0] mem_88_5_W0_addr;
  wire  mem_88_5_W0_clk;
  wire [7:0] mem_88_5_W0_data;
  wire  mem_88_5_W0_en;
  wire  mem_88_5_W0_mask;
  wire [25:0] mem_88_6_R0_addr;
  wire  mem_88_6_R0_clk;
  wire [7:0] mem_88_6_R0_data;
  wire  mem_88_6_R0_en;
  wire [25:0] mem_88_6_W0_addr;
  wire  mem_88_6_W0_clk;
  wire [7:0] mem_88_6_W0_data;
  wire  mem_88_6_W0_en;
  wire  mem_88_6_W0_mask;
  wire [25:0] mem_88_7_R0_addr;
  wire  mem_88_7_R0_clk;
  wire [7:0] mem_88_7_R0_data;
  wire  mem_88_7_R0_en;
  wire [25:0] mem_88_7_W0_addr;
  wire  mem_88_7_W0_clk;
  wire [7:0] mem_88_7_W0_data;
  wire  mem_88_7_W0_en;
  wire  mem_88_7_W0_mask;
  wire [25:0] mem_89_0_R0_addr;
  wire  mem_89_0_R0_clk;
  wire [7:0] mem_89_0_R0_data;
  wire  mem_89_0_R0_en;
  wire [25:0] mem_89_0_W0_addr;
  wire  mem_89_0_W0_clk;
  wire [7:0] mem_89_0_W0_data;
  wire  mem_89_0_W0_en;
  wire  mem_89_0_W0_mask;
  wire [25:0] mem_89_1_R0_addr;
  wire  mem_89_1_R0_clk;
  wire [7:0] mem_89_1_R0_data;
  wire  mem_89_1_R0_en;
  wire [25:0] mem_89_1_W0_addr;
  wire  mem_89_1_W0_clk;
  wire [7:0] mem_89_1_W0_data;
  wire  mem_89_1_W0_en;
  wire  mem_89_1_W0_mask;
  wire [25:0] mem_89_2_R0_addr;
  wire  mem_89_2_R0_clk;
  wire [7:0] mem_89_2_R0_data;
  wire  mem_89_2_R0_en;
  wire [25:0] mem_89_2_W0_addr;
  wire  mem_89_2_W0_clk;
  wire [7:0] mem_89_2_W0_data;
  wire  mem_89_2_W0_en;
  wire  mem_89_2_W0_mask;
  wire [25:0] mem_89_3_R0_addr;
  wire  mem_89_3_R0_clk;
  wire [7:0] mem_89_3_R0_data;
  wire  mem_89_3_R0_en;
  wire [25:0] mem_89_3_W0_addr;
  wire  mem_89_3_W0_clk;
  wire [7:0] mem_89_3_W0_data;
  wire  mem_89_3_W0_en;
  wire  mem_89_3_W0_mask;
  wire [25:0] mem_89_4_R0_addr;
  wire  mem_89_4_R0_clk;
  wire [7:0] mem_89_4_R0_data;
  wire  mem_89_4_R0_en;
  wire [25:0] mem_89_4_W0_addr;
  wire  mem_89_4_W0_clk;
  wire [7:0] mem_89_4_W0_data;
  wire  mem_89_4_W0_en;
  wire  mem_89_4_W0_mask;
  wire [25:0] mem_89_5_R0_addr;
  wire  mem_89_5_R0_clk;
  wire [7:0] mem_89_5_R0_data;
  wire  mem_89_5_R0_en;
  wire [25:0] mem_89_5_W0_addr;
  wire  mem_89_5_W0_clk;
  wire [7:0] mem_89_5_W0_data;
  wire  mem_89_5_W0_en;
  wire  mem_89_5_W0_mask;
  wire [25:0] mem_89_6_R0_addr;
  wire  mem_89_6_R0_clk;
  wire [7:0] mem_89_6_R0_data;
  wire  mem_89_6_R0_en;
  wire [25:0] mem_89_6_W0_addr;
  wire  mem_89_6_W0_clk;
  wire [7:0] mem_89_6_W0_data;
  wire  mem_89_6_W0_en;
  wire  mem_89_6_W0_mask;
  wire [25:0] mem_89_7_R0_addr;
  wire  mem_89_7_R0_clk;
  wire [7:0] mem_89_7_R0_data;
  wire  mem_89_7_R0_en;
  wire [25:0] mem_89_7_W0_addr;
  wire  mem_89_7_W0_clk;
  wire [7:0] mem_89_7_W0_data;
  wire  mem_89_7_W0_en;
  wire  mem_89_7_W0_mask;
  wire [25:0] mem_90_0_R0_addr;
  wire  mem_90_0_R0_clk;
  wire [7:0] mem_90_0_R0_data;
  wire  mem_90_0_R0_en;
  wire [25:0] mem_90_0_W0_addr;
  wire  mem_90_0_W0_clk;
  wire [7:0] mem_90_0_W0_data;
  wire  mem_90_0_W0_en;
  wire  mem_90_0_W0_mask;
  wire [25:0] mem_90_1_R0_addr;
  wire  mem_90_1_R0_clk;
  wire [7:0] mem_90_1_R0_data;
  wire  mem_90_1_R0_en;
  wire [25:0] mem_90_1_W0_addr;
  wire  mem_90_1_W0_clk;
  wire [7:0] mem_90_1_W0_data;
  wire  mem_90_1_W0_en;
  wire  mem_90_1_W0_mask;
  wire [25:0] mem_90_2_R0_addr;
  wire  mem_90_2_R0_clk;
  wire [7:0] mem_90_2_R0_data;
  wire  mem_90_2_R0_en;
  wire [25:0] mem_90_2_W0_addr;
  wire  mem_90_2_W0_clk;
  wire [7:0] mem_90_2_W0_data;
  wire  mem_90_2_W0_en;
  wire  mem_90_2_W0_mask;
  wire [25:0] mem_90_3_R0_addr;
  wire  mem_90_3_R0_clk;
  wire [7:0] mem_90_3_R0_data;
  wire  mem_90_3_R0_en;
  wire [25:0] mem_90_3_W0_addr;
  wire  mem_90_3_W0_clk;
  wire [7:0] mem_90_3_W0_data;
  wire  mem_90_3_W0_en;
  wire  mem_90_3_W0_mask;
  wire [25:0] mem_90_4_R0_addr;
  wire  mem_90_4_R0_clk;
  wire [7:0] mem_90_4_R0_data;
  wire  mem_90_4_R0_en;
  wire [25:0] mem_90_4_W0_addr;
  wire  mem_90_4_W0_clk;
  wire [7:0] mem_90_4_W0_data;
  wire  mem_90_4_W0_en;
  wire  mem_90_4_W0_mask;
  wire [25:0] mem_90_5_R0_addr;
  wire  mem_90_5_R0_clk;
  wire [7:0] mem_90_5_R0_data;
  wire  mem_90_5_R0_en;
  wire [25:0] mem_90_5_W0_addr;
  wire  mem_90_5_W0_clk;
  wire [7:0] mem_90_5_W0_data;
  wire  mem_90_5_W0_en;
  wire  mem_90_5_W0_mask;
  wire [25:0] mem_90_6_R0_addr;
  wire  mem_90_6_R0_clk;
  wire [7:0] mem_90_6_R0_data;
  wire  mem_90_6_R0_en;
  wire [25:0] mem_90_6_W0_addr;
  wire  mem_90_6_W0_clk;
  wire [7:0] mem_90_6_W0_data;
  wire  mem_90_6_W0_en;
  wire  mem_90_6_W0_mask;
  wire [25:0] mem_90_7_R0_addr;
  wire  mem_90_7_R0_clk;
  wire [7:0] mem_90_7_R0_data;
  wire  mem_90_7_R0_en;
  wire [25:0] mem_90_7_W0_addr;
  wire  mem_90_7_W0_clk;
  wire [7:0] mem_90_7_W0_data;
  wire  mem_90_7_W0_en;
  wire  mem_90_7_W0_mask;
  wire [25:0] mem_91_0_R0_addr;
  wire  mem_91_0_R0_clk;
  wire [7:0] mem_91_0_R0_data;
  wire  mem_91_0_R0_en;
  wire [25:0] mem_91_0_W0_addr;
  wire  mem_91_0_W0_clk;
  wire [7:0] mem_91_0_W0_data;
  wire  mem_91_0_W0_en;
  wire  mem_91_0_W0_mask;
  wire [25:0] mem_91_1_R0_addr;
  wire  mem_91_1_R0_clk;
  wire [7:0] mem_91_1_R0_data;
  wire  mem_91_1_R0_en;
  wire [25:0] mem_91_1_W0_addr;
  wire  mem_91_1_W0_clk;
  wire [7:0] mem_91_1_W0_data;
  wire  mem_91_1_W0_en;
  wire  mem_91_1_W0_mask;
  wire [25:0] mem_91_2_R0_addr;
  wire  mem_91_2_R0_clk;
  wire [7:0] mem_91_2_R0_data;
  wire  mem_91_2_R0_en;
  wire [25:0] mem_91_2_W0_addr;
  wire  mem_91_2_W0_clk;
  wire [7:0] mem_91_2_W0_data;
  wire  mem_91_2_W0_en;
  wire  mem_91_2_W0_mask;
  wire [25:0] mem_91_3_R0_addr;
  wire  mem_91_3_R0_clk;
  wire [7:0] mem_91_3_R0_data;
  wire  mem_91_3_R0_en;
  wire [25:0] mem_91_3_W0_addr;
  wire  mem_91_3_W0_clk;
  wire [7:0] mem_91_3_W0_data;
  wire  mem_91_3_W0_en;
  wire  mem_91_3_W0_mask;
  wire [25:0] mem_91_4_R0_addr;
  wire  mem_91_4_R0_clk;
  wire [7:0] mem_91_4_R0_data;
  wire  mem_91_4_R0_en;
  wire [25:0] mem_91_4_W0_addr;
  wire  mem_91_4_W0_clk;
  wire [7:0] mem_91_4_W0_data;
  wire  mem_91_4_W0_en;
  wire  mem_91_4_W0_mask;
  wire [25:0] mem_91_5_R0_addr;
  wire  mem_91_5_R0_clk;
  wire [7:0] mem_91_5_R0_data;
  wire  mem_91_5_R0_en;
  wire [25:0] mem_91_5_W0_addr;
  wire  mem_91_5_W0_clk;
  wire [7:0] mem_91_5_W0_data;
  wire  mem_91_5_W0_en;
  wire  mem_91_5_W0_mask;
  wire [25:0] mem_91_6_R0_addr;
  wire  mem_91_6_R0_clk;
  wire [7:0] mem_91_6_R0_data;
  wire  mem_91_6_R0_en;
  wire [25:0] mem_91_6_W0_addr;
  wire  mem_91_6_W0_clk;
  wire [7:0] mem_91_6_W0_data;
  wire  mem_91_6_W0_en;
  wire  mem_91_6_W0_mask;
  wire [25:0] mem_91_7_R0_addr;
  wire  mem_91_7_R0_clk;
  wire [7:0] mem_91_7_R0_data;
  wire  mem_91_7_R0_en;
  wire [25:0] mem_91_7_W0_addr;
  wire  mem_91_7_W0_clk;
  wire [7:0] mem_91_7_W0_data;
  wire  mem_91_7_W0_en;
  wire  mem_91_7_W0_mask;
  wire [25:0] mem_92_0_R0_addr;
  wire  mem_92_0_R0_clk;
  wire [7:0] mem_92_0_R0_data;
  wire  mem_92_0_R0_en;
  wire [25:0] mem_92_0_W0_addr;
  wire  mem_92_0_W0_clk;
  wire [7:0] mem_92_0_W0_data;
  wire  mem_92_0_W0_en;
  wire  mem_92_0_W0_mask;
  wire [25:0] mem_92_1_R0_addr;
  wire  mem_92_1_R0_clk;
  wire [7:0] mem_92_1_R0_data;
  wire  mem_92_1_R0_en;
  wire [25:0] mem_92_1_W0_addr;
  wire  mem_92_1_W0_clk;
  wire [7:0] mem_92_1_W0_data;
  wire  mem_92_1_W0_en;
  wire  mem_92_1_W0_mask;
  wire [25:0] mem_92_2_R0_addr;
  wire  mem_92_2_R0_clk;
  wire [7:0] mem_92_2_R0_data;
  wire  mem_92_2_R0_en;
  wire [25:0] mem_92_2_W0_addr;
  wire  mem_92_2_W0_clk;
  wire [7:0] mem_92_2_W0_data;
  wire  mem_92_2_W0_en;
  wire  mem_92_2_W0_mask;
  wire [25:0] mem_92_3_R0_addr;
  wire  mem_92_3_R0_clk;
  wire [7:0] mem_92_3_R0_data;
  wire  mem_92_3_R0_en;
  wire [25:0] mem_92_3_W0_addr;
  wire  mem_92_3_W0_clk;
  wire [7:0] mem_92_3_W0_data;
  wire  mem_92_3_W0_en;
  wire  mem_92_3_W0_mask;
  wire [25:0] mem_92_4_R0_addr;
  wire  mem_92_4_R0_clk;
  wire [7:0] mem_92_4_R0_data;
  wire  mem_92_4_R0_en;
  wire [25:0] mem_92_4_W0_addr;
  wire  mem_92_4_W0_clk;
  wire [7:0] mem_92_4_W0_data;
  wire  mem_92_4_W0_en;
  wire  mem_92_4_W0_mask;
  wire [25:0] mem_92_5_R0_addr;
  wire  mem_92_5_R0_clk;
  wire [7:0] mem_92_5_R0_data;
  wire  mem_92_5_R0_en;
  wire [25:0] mem_92_5_W0_addr;
  wire  mem_92_5_W0_clk;
  wire [7:0] mem_92_5_W0_data;
  wire  mem_92_5_W0_en;
  wire  mem_92_5_W0_mask;
  wire [25:0] mem_92_6_R0_addr;
  wire  mem_92_6_R0_clk;
  wire [7:0] mem_92_6_R0_data;
  wire  mem_92_6_R0_en;
  wire [25:0] mem_92_6_W0_addr;
  wire  mem_92_6_W0_clk;
  wire [7:0] mem_92_6_W0_data;
  wire  mem_92_6_W0_en;
  wire  mem_92_6_W0_mask;
  wire [25:0] mem_92_7_R0_addr;
  wire  mem_92_7_R0_clk;
  wire [7:0] mem_92_7_R0_data;
  wire  mem_92_7_R0_en;
  wire [25:0] mem_92_7_W0_addr;
  wire  mem_92_7_W0_clk;
  wire [7:0] mem_92_7_W0_data;
  wire  mem_92_7_W0_en;
  wire  mem_92_7_W0_mask;
  wire [25:0] mem_93_0_R0_addr;
  wire  mem_93_0_R0_clk;
  wire [7:0] mem_93_0_R0_data;
  wire  mem_93_0_R0_en;
  wire [25:0] mem_93_0_W0_addr;
  wire  mem_93_0_W0_clk;
  wire [7:0] mem_93_0_W0_data;
  wire  mem_93_0_W0_en;
  wire  mem_93_0_W0_mask;
  wire [25:0] mem_93_1_R0_addr;
  wire  mem_93_1_R0_clk;
  wire [7:0] mem_93_1_R0_data;
  wire  mem_93_1_R0_en;
  wire [25:0] mem_93_1_W0_addr;
  wire  mem_93_1_W0_clk;
  wire [7:0] mem_93_1_W0_data;
  wire  mem_93_1_W0_en;
  wire  mem_93_1_W0_mask;
  wire [25:0] mem_93_2_R0_addr;
  wire  mem_93_2_R0_clk;
  wire [7:0] mem_93_2_R0_data;
  wire  mem_93_2_R0_en;
  wire [25:0] mem_93_2_W0_addr;
  wire  mem_93_2_W0_clk;
  wire [7:0] mem_93_2_W0_data;
  wire  mem_93_2_W0_en;
  wire  mem_93_2_W0_mask;
  wire [25:0] mem_93_3_R0_addr;
  wire  mem_93_3_R0_clk;
  wire [7:0] mem_93_3_R0_data;
  wire  mem_93_3_R0_en;
  wire [25:0] mem_93_3_W0_addr;
  wire  mem_93_3_W0_clk;
  wire [7:0] mem_93_3_W0_data;
  wire  mem_93_3_W0_en;
  wire  mem_93_3_W0_mask;
  wire [25:0] mem_93_4_R0_addr;
  wire  mem_93_4_R0_clk;
  wire [7:0] mem_93_4_R0_data;
  wire  mem_93_4_R0_en;
  wire [25:0] mem_93_4_W0_addr;
  wire  mem_93_4_W0_clk;
  wire [7:0] mem_93_4_W0_data;
  wire  mem_93_4_W0_en;
  wire  mem_93_4_W0_mask;
  wire [25:0] mem_93_5_R0_addr;
  wire  mem_93_5_R0_clk;
  wire [7:0] mem_93_5_R0_data;
  wire  mem_93_5_R0_en;
  wire [25:0] mem_93_5_W0_addr;
  wire  mem_93_5_W0_clk;
  wire [7:0] mem_93_5_W0_data;
  wire  mem_93_5_W0_en;
  wire  mem_93_5_W0_mask;
  wire [25:0] mem_93_6_R0_addr;
  wire  mem_93_6_R0_clk;
  wire [7:0] mem_93_6_R0_data;
  wire  mem_93_6_R0_en;
  wire [25:0] mem_93_6_W0_addr;
  wire  mem_93_6_W0_clk;
  wire [7:0] mem_93_6_W0_data;
  wire  mem_93_6_W0_en;
  wire  mem_93_6_W0_mask;
  wire [25:0] mem_93_7_R0_addr;
  wire  mem_93_7_R0_clk;
  wire [7:0] mem_93_7_R0_data;
  wire  mem_93_7_R0_en;
  wire [25:0] mem_93_7_W0_addr;
  wire  mem_93_7_W0_clk;
  wire [7:0] mem_93_7_W0_data;
  wire  mem_93_7_W0_en;
  wire  mem_93_7_W0_mask;
  wire [25:0] mem_94_0_R0_addr;
  wire  mem_94_0_R0_clk;
  wire [7:0] mem_94_0_R0_data;
  wire  mem_94_0_R0_en;
  wire [25:0] mem_94_0_W0_addr;
  wire  mem_94_0_W0_clk;
  wire [7:0] mem_94_0_W0_data;
  wire  mem_94_0_W0_en;
  wire  mem_94_0_W0_mask;
  wire [25:0] mem_94_1_R0_addr;
  wire  mem_94_1_R0_clk;
  wire [7:0] mem_94_1_R0_data;
  wire  mem_94_1_R0_en;
  wire [25:0] mem_94_1_W0_addr;
  wire  mem_94_1_W0_clk;
  wire [7:0] mem_94_1_W0_data;
  wire  mem_94_1_W0_en;
  wire  mem_94_1_W0_mask;
  wire [25:0] mem_94_2_R0_addr;
  wire  mem_94_2_R0_clk;
  wire [7:0] mem_94_2_R0_data;
  wire  mem_94_2_R0_en;
  wire [25:0] mem_94_2_W0_addr;
  wire  mem_94_2_W0_clk;
  wire [7:0] mem_94_2_W0_data;
  wire  mem_94_2_W0_en;
  wire  mem_94_2_W0_mask;
  wire [25:0] mem_94_3_R0_addr;
  wire  mem_94_3_R0_clk;
  wire [7:0] mem_94_3_R0_data;
  wire  mem_94_3_R0_en;
  wire [25:0] mem_94_3_W0_addr;
  wire  mem_94_3_W0_clk;
  wire [7:0] mem_94_3_W0_data;
  wire  mem_94_3_W0_en;
  wire  mem_94_3_W0_mask;
  wire [25:0] mem_94_4_R0_addr;
  wire  mem_94_4_R0_clk;
  wire [7:0] mem_94_4_R0_data;
  wire  mem_94_4_R0_en;
  wire [25:0] mem_94_4_W0_addr;
  wire  mem_94_4_W0_clk;
  wire [7:0] mem_94_4_W0_data;
  wire  mem_94_4_W0_en;
  wire  mem_94_4_W0_mask;
  wire [25:0] mem_94_5_R0_addr;
  wire  mem_94_5_R0_clk;
  wire [7:0] mem_94_5_R0_data;
  wire  mem_94_5_R0_en;
  wire [25:0] mem_94_5_W0_addr;
  wire  mem_94_5_W0_clk;
  wire [7:0] mem_94_5_W0_data;
  wire  mem_94_5_W0_en;
  wire  mem_94_5_W0_mask;
  wire [25:0] mem_94_6_R0_addr;
  wire  mem_94_6_R0_clk;
  wire [7:0] mem_94_6_R0_data;
  wire  mem_94_6_R0_en;
  wire [25:0] mem_94_6_W0_addr;
  wire  mem_94_6_W0_clk;
  wire [7:0] mem_94_6_W0_data;
  wire  mem_94_6_W0_en;
  wire  mem_94_6_W0_mask;
  wire [25:0] mem_94_7_R0_addr;
  wire  mem_94_7_R0_clk;
  wire [7:0] mem_94_7_R0_data;
  wire  mem_94_7_R0_en;
  wire [25:0] mem_94_7_W0_addr;
  wire  mem_94_7_W0_clk;
  wire [7:0] mem_94_7_W0_data;
  wire  mem_94_7_W0_en;
  wire  mem_94_7_W0_mask;
  wire [25:0] mem_95_0_R0_addr;
  wire  mem_95_0_R0_clk;
  wire [7:0] mem_95_0_R0_data;
  wire  mem_95_0_R0_en;
  wire [25:0] mem_95_0_W0_addr;
  wire  mem_95_0_W0_clk;
  wire [7:0] mem_95_0_W0_data;
  wire  mem_95_0_W0_en;
  wire  mem_95_0_W0_mask;
  wire [25:0] mem_95_1_R0_addr;
  wire  mem_95_1_R0_clk;
  wire [7:0] mem_95_1_R0_data;
  wire  mem_95_1_R0_en;
  wire [25:0] mem_95_1_W0_addr;
  wire  mem_95_1_W0_clk;
  wire [7:0] mem_95_1_W0_data;
  wire  mem_95_1_W0_en;
  wire  mem_95_1_W0_mask;
  wire [25:0] mem_95_2_R0_addr;
  wire  mem_95_2_R0_clk;
  wire [7:0] mem_95_2_R0_data;
  wire  mem_95_2_R0_en;
  wire [25:0] mem_95_2_W0_addr;
  wire  mem_95_2_W0_clk;
  wire [7:0] mem_95_2_W0_data;
  wire  mem_95_2_W0_en;
  wire  mem_95_2_W0_mask;
  wire [25:0] mem_95_3_R0_addr;
  wire  mem_95_3_R0_clk;
  wire [7:0] mem_95_3_R0_data;
  wire  mem_95_3_R0_en;
  wire [25:0] mem_95_3_W0_addr;
  wire  mem_95_3_W0_clk;
  wire [7:0] mem_95_3_W0_data;
  wire  mem_95_3_W0_en;
  wire  mem_95_3_W0_mask;
  wire [25:0] mem_95_4_R0_addr;
  wire  mem_95_4_R0_clk;
  wire [7:0] mem_95_4_R0_data;
  wire  mem_95_4_R0_en;
  wire [25:0] mem_95_4_W0_addr;
  wire  mem_95_4_W0_clk;
  wire [7:0] mem_95_4_W0_data;
  wire  mem_95_4_W0_en;
  wire  mem_95_4_W0_mask;
  wire [25:0] mem_95_5_R0_addr;
  wire  mem_95_5_R0_clk;
  wire [7:0] mem_95_5_R0_data;
  wire  mem_95_5_R0_en;
  wire [25:0] mem_95_5_W0_addr;
  wire  mem_95_5_W0_clk;
  wire [7:0] mem_95_5_W0_data;
  wire  mem_95_5_W0_en;
  wire  mem_95_5_W0_mask;
  wire [25:0] mem_95_6_R0_addr;
  wire  mem_95_6_R0_clk;
  wire [7:0] mem_95_6_R0_data;
  wire  mem_95_6_R0_en;
  wire [25:0] mem_95_6_W0_addr;
  wire  mem_95_6_W0_clk;
  wire [7:0] mem_95_6_W0_data;
  wire  mem_95_6_W0_en;
  wire  mem_95_6_W0_mask;
  wire [25:0] mem_95_7_R0_addr;
  wire  mem_95_7_R0_clk;
  wire [7:0] mem_95_7_R0_data;
  wire  mem_95_7_R0_en;
  wire [25:0] mem_95_7_W0_addr;
  wire  mem_95_7_W0_clk;
  wire [7:0] mem_95_7_W0_data;
  wire  mem_95_7_W0_en;
  wire  mem_95_7_W0_mask;
  wire [25:0] mem_96_0_R0_addr;
  wire  mem_96_0_R0_clk;
  wire [7:0] mem_96_0_R0_data;
  wire  mem_96_0_R0_en;
  wire [25:0] mem_96_0_W0_addr;
  wire  mem_96_0_W0_clk;
  wire [7:0] mem_96_0_W0_data;
  wire  mem_96_0_W0_en;
  wire  mem_96_0_W0_mask;
  wire [25:0] mem_96_1_R0_addr;
  wire  mem_96_1_R0_clk;
  wire [7:0] mem_96_1_R0_data;
  wire  mem_96_1_R0_en;
  wire [25:0] mem_96_1_W0_addr;
  wire  mem_96_1_W0_clk;
  wire [7:0] mem_96_1_W0_data;
  wire  mem_96_1_W0_en;
  wire  mem_96_1_W0_mask;
  wire [25:0] mem_96_2_R0_addr;
  wire  mem_96_2_R0_clk;
  wire [7:0] mem_96_2_R0_data;
  wire  mem_96_2_R0_en;
  wire [25:0] mem_96_2_W0_addr;
  wire  mem_96_2_W0_clk;
  wire [7:0] mem_96_2_W0_data;
  wire  mem_96_2_W0_en;
  wire  mem_96_2_W0_mask;
  wire [25:0] mem_96_3_R0_addr;
  wire  mem_96_3_R0_clk;
  wire [7:0] mem_96_3_R0_data;
  wire  mem_96_3_R0_en;
  wire [25:0] mem_96_3_W0_addr;
  wire  mem_96_3_W0_clk;
  wire [7:0] mem_96_3_W0_data;
  wire  mem_96_3_W0_en;
  wire  mem_96_3_W0_mask;
  wire [25:0] mem_96_4_R0_addr;
  wire  mem_96_4_R0_clk;
  wire [7:0] mem_96_4_R0_data;
  wire  mem_96_4_R0_en;
  wire [25:0] mem_96_4_W0_addr;
  wire  mem_96_4_W0_clk;
  wire [7:0] mem_96_4_W0_data;
  wire  mem_96_4_W0_en;
  wire  mem_96_4_W0_mask;
  wire [25:0] mem_96_5_R0_addr;
  wire  mem_96_5_R0_clk;
  wire [7:0] mem_96_5_R0_data;
  wire  mem_96_5_R0_en;
  wire [25:0] mem_96_5_W0_addr;
  wire  mem_96_5_W0_clk;
  wire [7:0] mem_96_5_W0_data;
  wire  mem_96_5_W0_en;
  wire  mem_96_5_W0_mask;
  wire [25:0] mem_96_6_R0_addr;
  wire  mem_96_6_R0_clk;
  wire [7:0] mem_96_6_R0_data;
  wire  mem_96_6_R0_en;
  wire [25:0] mem_96_6_W0_addr;
  wire  mem_96_6_W0_clk;
  wire [7:0] mem_96_6_W0_data;
  wire  mem_96_6_W0_en;
  wire  mem_96_6_W0_mask;
  wire [25:0] mem_96_7_R0_addr;
  wire  mem_96_7_R0_clk;
  wire [7:0] mem_96_7_R0_data;
  wire  mem_96_7_R0_en;
  wire [25:0] mem_96_7_W0_addr;
  wire  mem_96_7_W0_clk;
  wire [7:0] mem_96_7_W0_data;
  wire  mem_96_7_W0_en;
  wire  mem_96_7_W0_mask;
  wire [25:0] mem_97_0_R0_addr;
  wire  mem_97_0_R0_clk;
  wire [7:0] mem_97_0_R0_data;
  wire  mem_97_0_R0_en;
  wire [25:0] mem_97_0_W0_addr;
  wire  mem_97_0_W0_clk;
  wire [7:0] mem_97_0_W0_data;
  wire  mem_97_0_W0_en;
  wire  mem_97_0_W0_mask;
  wire [25:0] mem_97_1_R0_addr;
  wire  mem_97_1_R0_clk;
  wire [7:0] mem_97_1_R0_data;
  wire  mem_97_1_R0_en;
  wire [25:0] mem_97_1_W0_addr;
  wire  mem_97_1_W0_clk;
  wire [7:0] mem_97_1_W0_data;
  wire  mem_97_1_W0_en;
  wire  mem_97_1_W0_mask;
  wire [25:0] mem_97_2_R0_addr;
  wire  mem_97_2_R0_clk;
  wire [7:0] mem_97_2_R0_data;
  wire  mem_97_2_R0_en;
  wire [25:0] mem_97_2_W0_addr;
  wire  mem_97_2_W0_clk;
  wire [7:0] mem_97_2_W0_data;
  wire  mem_97_2_W0_en;
  wire  mem_97_2_W0_mask;
  wire [25:0] mem_97_3_R0_addr;
  wire  mem_97_3_R0_clk;
  wire [7:0] mem_97_3_R0_data;
  wire  mem_97_3_R0_en;
  wire [25:0] mem_97_3_W0_addr;
  wire  mem_97_3_W0_clk;
  wire [7:0] mem_97_3_W0_data;
  wire  mem_97_3_W0_en;
  wire  mem_97_3_W0_mask;
  wire [25:0] mem_97_4_R0_addr;
  wire  mem_97_4_R0_clk;
  wire [7:0] mem_97_4_R0_data;
  wire  mem_97_4_R0_en;
  wire [25:0] mem_97_4_W0_addr;
  wire  mem_97_4_W0_clk;
  wire [7:0] mem_97_4_W0_data;
  wire  mem_97_4_W0_en;
  wire  mem_97_4_W0_mask;
  wire [25:0] mem_97_5_R0_addr;
  wire  mem_97_5_R0_clk;
  wire [7:0] mem_97_5_R0_data;
  wire  mem_97_5_R0_en;
  wire [25:0] mem_97_5_W0_addr;
  wire  mem_97_5_W0_clk;
  wire [7:0] mem_97_5_W0_data;
  wire  mem_97_5_W0_en;
  wire  mem_97_5_W0_mask;
  wire [25:0] mem_97_6_R0_addr;
  wire  mem_97_6_R0_clk;
  wire [7:0] mem_97_6_R0_data;
  wire  mem_97_6_R0_en;
  wire [25:0] mem_97_6_W0_addr;
  wire  mem_97_6_W0_clk;
  wire [7:0] mem_97_6_W0_data;
  wire  mem_97_6_W0_en;
  wire  mem_97_6_W0_mask;
  wire [25:0] mem_97_7_R0_addr;
  wire  mem_97_7_R0_clk;
  wire [7:0] mem_97_7_R0_data;
  wire  mem_97_7_R0_en;
  wire [25:0] mem_97_7_W0_addr;
  wire  mem_97_7_W0_clk;
  wire [7:0] mem_97_7_W0_data;
  wire  mem_97_7_W0_en;
  wire  mem_97_7_W0_mask;
  wire [25:0] mem_98_0_R0_addr;
  wire  mem_98_0_R0_clk;
  wire [7:0] mem_98_0_R0_data;
  wire  mem_98_0_R0_en;
  wire [25:0] mem_98_0_W0_addr;
  wire  mem_98_0_W0_clk;
  wire [7:0] mem_98_0_W0_data;
  wire  mem_98_0_W0_en;
  wire  mem_98_0_W0_mask;
  wire [25:0] mem_98_1_R0_addr;
  wire  mem_98_1_R0_clk;
  wire [7:0] mem_98_1_R0_data;
  wire  mem_98_1_R0_en;
  wire [25:0] mem_98_1_W0_addr;
  wire  mem_98_1_W0_clk;
  wire [7:0] mem_98_1_W0_data;
  wire  mem_98_1_W0_en;
  wire  mem_98_1_W0_mask;
  wire [25:0] mem_98_2_R0_addr;
  wire  mem_98_2_R0_clk;
  wire [7:0] mem_98_2_R0_data;
  wire  mem_98_2_R0_en;
  wire [25:0] mem_98_2_W0_addr;
  wire  mem_98_2_W0_clk;
  wire [7:0] mem_98_2_W0_data;
  wire  mem_98_2_W0_en;
  wire  mem_98_2_W0_mask;
  wire [25:0] mem_98_3_R0_addr;
  wire  mem_98_3_R0_clk;
  wire [7:0] mem_98_3_R0_data;
  wire  mem_98_3_R0_en;
  wire [25:0] mem_98_3_W0_addr;
  wire  mem_98_3_W0_clk;
  wire [7:0] mem_98_3_W0_data;
  wire  mem_98_3_W0_en;
  wire  mem_98_3_W0_mask;
  wire [25:0] mem_98_4_R0_addr;
  wire  mem_98_4_R0_clk;
  wire [7:0] mem_98_4_R0_data;
  wire  mem_98_4_R0_en;
  wire [25:0] mem_98_4_W0_addr;
  wire  mem_98_4_W0_clk;
  wire [7:0] mem_98_4_W0_data;
  wire  mem_98_4_W0_en;
  wire  mem_98_4_W0_mask;
  wire [25:0] mem_98_5_R0_addr;
  wire  mem_98_5_R0_clk;
  wire [7:0] mem_98_5_R0_data;
  wire  mem_98_5_R0_en;
  wire [25:0] mem_98_5_W0_addr;
  wire  mem_98_5_W0_clk;
  wire [7:0] mem_98_5_W0_data;
  wire  mem_98_5_W0_en;
  wire  mem_98_5_W0_mask;
  wire [25:0] mem_98_6_R0_addr;
  wire  mem_98_6_R0_clk;
  wire [7:0] mem_98_6_R0_data;
  wire  mem_98_6_R0_en;
  wire [25:0] mem_98_6_W0_addr;
  wire  mem_98_6_W0_clk;
  wire [7:0] mem_98_6_W0_data;
  wire  mem_98_6_W0_en;
  wire  mem_98_6_W0_mask;
  wire [25:0] mem_98_7_R0_addr;
  wire  mem_98_7_R0_clk;
  wire [7:0] mem_98_7_R0_data;
  wire  mem_98_7_R0_en;
  wire [25:0] mem_98_7_W0_addr;
  wire  mem_98_7_W0_clk;
  wire [7:0] mem_98_7_W0_data;
  wire  mem_98_7_W0_en;
  wire  mem_98_7_W0_mask;
  wire [25:0] mem_99_0_R0_addr;
  wire  mem_99_0_R0_clk;
  wire [7:0] mem_99_0_R0_data;
  wire  mem_99_0_R0_en;
  wire [25:0] mem_99_0_W0_addr;
  wire  mem_99_0_W0_clk;
  wire [7:0] mem_99_0_W0_data;
  wire  mem_99_0_W0_en;
  wire  mem_99_0_W0_mask;
  wire [25:0] mem_99_1_R0_addr;
  wire  mem_99_1_R0_clk;
  wire [7:0] mem_99_1_R0_data;
  wire  mem_99_1_R0_en;
  wire [25:0] mem_99_1_W0_addr;
  wire  mem_99_1_W0_clk;
  wire [7:0] mem_99_1_W0_data;
  wire  mem_99_1_W0_en;
  wire  mem_99_1_W0_mask;
  wire [25:0] mem_99_2_R0_addr;
  wire  mem_99_2_R0_clk;
  wire [7:0] mem_99_2_R0_data;
  wire  mem_99_2_R0_en;
  wire [25:0] mem_99_2_W0_addr;
  wire  mem_99_2_W0_clk;
  wire [7:0] mem_99_2_W0_data;
  wire  mem_99_2_W0_en;
  wire  mem_99_2_W0_mask;
  wire [25:0] mem_99_3_R0_addr;
  wire  mem_99_3_R0_clk;
  wire [7:0] mem_99_3_R0_data;
  wire  mem_99_3_R0_en;
  wire [25:0] mem_99_3_W0_addr;
  wire  mem_99_3_W0_clk;
  wire [7:0] mem_99_3_W0_data;
  wire  mem_99_3_W0_en;
  wire  mem_99_3_W0_mask;
  wire [25:0] mem_99_4_R0_addr;
  wire  mem_99_4_R0_clk;
  wire [7:0] mem_99_4_R0_data;
  wire  mem_99_4_R0_en;
  wire [25:0] mem_99_4_W0_addr;
  wire  mem_99_4_W0_clk;
  wire [7:0] mem_99_4_W0_data;
  wire  mem_99_4_W0_en;
  wire  mem_99_4_W0_mask;
  wire [25:0] mem_99_5_R0_addr;
  wire  mem_99_5_R0_clk;
  wire [7:0] mem_99_5_R0_data;
  wire  mem_99_5_R0_en;
  wire [25:0] mem_99_5_W0_addr;
  wire  mem_99_5_W0_clk;
  wire [7:0] mem_99_5_W0_data;
  wire  mem_99_5_W0_en;
  wire  mem_99_5_W0_mask;
  wire [25:0] mem_99_6_R0_addr;
  wire  mem_99_6_R0_clk;
  wire [7:0] mem_99_6_R0_data;
  wire  mem_99_6_R0_en;
  wire [25:0] mem_99_6_W0_addr;
  wire  mem_99_6_W0_clk;
  wire [7:0] mem_99_6_W0_data;
  wire  mem_99_6_W0_en;
  wire  mem_99_6_W0_mask;
  wire [25:0] mem_99_7_R0_addr;
  wire  mem_99_7_R0_clk;
  wire [7:0] mem_99_7_R0_data;
  wire  mem_99_7_R0_en;
  wire [25:0] mem_99_7_W0_addr;
  wire  mem_99_7_W0_clk;
  wire [7:0] mem_99_7_W0_data;
  wire  mem_99_7_W0_en;
  wire  mem_99_7_W0_mask;
  wire [25:0] mem_100_0_R0_addr;
  wire  mem_100_0_R0_clk;
  wire [7:0] mem_100_0_R0_data;
  wire  mem_100_0_R0_en;
  wire [25:0] mem_100_0_W0_addr;
  wire  mem_100_0_W0_clk;
  wire [7:0] mem_100_0_W0_data;
  wire  mem_100_0_W0_en;
  wire  mem_100_0_W0_mask;
  wire [25:0] mem_100_1_R0_addr;
  wire  mem_100_1_R0_clk;
  wire [7:0] mem_100_1_R0_data;
  wire  mem_100_1_R0_en;
  wire [25:0] mem_100_1_W0_addr;
  wire  mem_100_1_W0_clk;
  wire [7:0] mem_100_1_W0_data;
  wire  mem_100_1_W0_en;
  wire  mem_100_1_W0_mask;
  wire [25:0] mem_100_2_R0_addr;
  wire  mem_100_2_R0_clk;
  wire [7:0] mem_100_2_R0_data;
  wire  mem_100_2_R0_en;
  wire [25:0] mem_100_2_W0_addr;
  wire  mem_100_2_W0_clk;
  wire [7:0] mem_100_2_W0_data;
  wire  mem_100_2_W0_en;
  wire  mem_100_2_W0_mask;
  wire [25:0] mem_100_3_R0_addr;
  wire  mem_100_3_R0_clk;
  wire [7:0] mem_100_3_R0_data;
  wire  mem_100_3_R0_en;
  wire [25:0] mem_100_3_W0_addr;
  wire  mem_100_3_W0_clk;
  wire [7:0] mem_100_3_W0_data;
  wire  mem_100_3_W0_en;
  wire  mem_100_3_W0_mask;
  wire [25:0] mem_100_4_R0_addr;
  wire  mem_100_4_R0_clk;
  wire [7:0] mem_100_4_R0_data;
  wire  mem_100_4_R0_en;
  wire [25:0] mem_100_4_W0_addr;
  wire  mem_100_4_W0_clk;
  wire [7:0] mem_100_4_W0_data;
  wire  mem_100_4_W0_en;
  wire  mem_100_4_W0_mask;
  wire [25:0] mem_100_5_R0_addr;
  wire  mem_100_5_R0_clk;
  wire [7:0] mem_100_5_R0_data;
  wire  mem_100_5_R0_en;
  wire [25:0] mem_100_5_W0_addr;
  wire  mem_100_5_W0_clk;
  wire [7:0] mem_100_5_W0_data;
  wire  mem_100_5_W0_en;
  wire  mem_100_5_W0_mask;
  wire [25:0] mem_100_6_R0_addr;
  wire  mem_100_6_R0_clk;
  wire [7:0] mem_100_6_R0_data;
  wire  mem_100_6_R0_en;
  wire [25:0] mem_100_6_W0_addr;
  wire  mem_100_6_W0_clk;
  wire [7:0] mem_100_6_W0_data;
  wire  mem_100_6_W0_en;
  wire  mem_100_6_W0_mask;
  wire [25:0] mem_100_7_R0_addr;
  wire  mem_100_7_R0_clk;
  wire [7:0] mem_100_7_R0_data;
  wire  mem_100_7_R0_en;
  wire [25:0] mem_100_7_W0_addr;
  wire  mem_100_7_W0_clk;
  wire [7:0] mem_100_7_W0_data;
  wire  mem_100_7_W0_en;
  wire  mem_100_7_W0_mask;
  wire [25:0] mem_101_0_R0_addr;
  wire  mem_101_0_R0_clk;
  wire [7:0] mem_101_0_R0_data;
  wire  mem_101_0_R0_en;
  wire [25:0] mem_101_0_W0_addr;
  wire  mem_101_0_W0_clk;
  wire [7:0] mem_101_0_W0_data;
  wire  mem_101_0_W0_en;
  wire  mem_101_0_W0_mask;
  wire [25:0] mem_101_1_R0_addr;
  wire  mem_101_1_R0_clk;
  wire [7:0] mem_101_1_R0_data;
  wire  mem_101_1_R0_en;
  wire [25:0] mem_101_1_W0_addr;
  wire  mem_101_1_W0_clk;
  wire [7:0] mem_101_1_W0_data;
  wire  mem_101_1_W0_en;
  wire  mem_101_1_W0_mask;
  wire [25:0] mem_101_2_R0_addr;
  wire  mem_101_2_R0_clk;
  wire [7:0] mem_101_2_R0_data;
  wire  mem_101_2_R0_en;
  wire [25:0] mem_101_2_W0_addr;
  wire  mem_101_2_W0_clk;
  wire [7:0] mem_101_2_W0_data;
  wire  mem_101_2_W0_en;
  wire  mem_101_2_W0_mask;
  wire [25:0] mem_101_3_R0_addr;
  wire  mem_101_3_R0_clk;
  wire [7:0] mem_101_3_R0_data;
  wire  mem_101_3_R0_en;
  wire [25:0] mem_101_3_W0_addr;
  wire  mem_101_3_W0_clk;
  wire [7:0] mem_101_3_W0_data;
  wire  mem_101_3_W0_en;
  wire  mem_101_3_W0_mask;
  wire [25:0] mem_101_4_R0_addr;
  wire  mem_101_4_R0_clk;
  wire [7:0] mem_101_4_R0_data;
  wire  mem_101_4_R0_en;
  wire [25:0] mem_101_4_W0_addr;
  wire  mem_101_4_W0_clk;
  wire [7:0] mem_101_4_W0_data;
  wire  mem_101_4_W0_en;
  wire  mem_101_4_W0_mask;
  wire [25:0] mem_101_5_R0_addr;
  wire  mem_101_5_R0_clk;
  wire [7:0] mem_101_5_R0_data;
  wire  mem_101_5_R0_en;
  wire [25:0] mem_101_5_W0_addr;
  wire  mem_101_5_W0_clk;
  wire [7:0] mem_101_5_W0_data;
  wire  mem_101_5_W0_en;
  wire  mem_101_5_W0_mask;
  wire [25:0] mem_101_6_R0_addr;
  wire  mem_101_6_R0_clk;
  wire [7:0] mem_101_6_R0_data;
  wire  mem_101_6_R0_en;
  wire [25:0] mem_101_6_W0_addr;
  wire  mem_101_6_W0_clk;
  wire [7:0] mem_101_6_W0_data;
  wire  mem_101_6_W0_en;
  wire  mem_101_6_W0_mask;
  wire [25:0] mem_101_7_R0_addr;
  wire  mem_101_7_R0_clk;
  wire [7:0] mem_101_7_R0_data;
  wire  mem_101_7_R0_en;
  wire [25:0] mem_101_7_W0_addr;
  wire  mem_101_7_W0_clk;
  wire [7:0] mem_101_7_W0_data;
  wire  mem_101_7_W0_en;
  wire  mem_101_7_W0_mask;
  wire [25:0] mem_102_0_R0_addr;
  wire  mem_102_0_R0_clk;
  wire [7:0] mem_102_0_R0_data;
  wire  mem_102_0_R0_en;
  wire [25:0] mem_102_0_W0_addr;
  wire  mem_102_0_W0_clk;
  wire [7:0] mem_102_0_W0_data;
  wire  mem_102_0_W0_en;
  wire  mem_102_0_W0_mask;
  wire [25:0] mem_102_1_R0_addr;
  wire  mem_102_1_R0_clk;
  wire [7:0] mem_102_1_R0_data;
  wire  mem_102_1_R0_en;
  wire [25:0] mem_102_1_W0_addr;
  wire  mem_102_1_W0_clk;
  wire [7:0] mem_102_1_W0_data;
  wire  mem_102_1_W0_en;
  wire  mem_102_1_W0_mask;
  wire [25:0] mem_102_2_R0_addr;
  wire  mem_102_2_R0_clk;
  wire [7:0] mem_102_2_R0_data;
  wire  mem_102_2_R0_en;
  wire [25:0] mem_102_2_W0_addr;
  wire  mem_102_2_W0_clk;
  wire [7:0] mem_102_2_W0_data;
  wire  mem_102_2_W0_en;
  wire  mem_102_2_W0_mask;
  wire [25:0] mem_102_3_R0_addr;
  wire  mem_102_3_R0_clk;
  wire [7:0] mem_102_3_R0_data;
  wire  mem_102_3_R0_en;
  wire [25:0] mem_102_3_W0_addr;
  wire  mem_102_3_W0_clk;
  wire [7:0] mem_102_3_W0_data;
  wire  mem_102_3_W0_en;
  wire  mem_102_3_W0_mask;
  wire [25:0] mem_102_4_R0_addr;
  wire  mem_102_4_R0_clk;
  wire [7:0] mem_102_4_R0_data;
  wire  mem_102_4_R0_en;
  wire [25:0] mem_102_4_W0_addr;
  wire  mem_102_4_W0_clk;
  wire [7:0] mem_102_4_W0_data;
  wire  mem_102_4_W0_en;
  wire  mem_102_4_W0_mask;
  wire [25:0] mem_102_5_R0_addr;
  wire  mem_102_5_R0_clk;
  wire [7:0] mem_102_5_R0_data;
  wire  mem_102_5_R0_en;
  wire [25:0] mem_102_5_W0_addr;
  wire  mem_102_5_W0_clk;
  wire [7:0] mem_102_5_W0_data;
  wire  mem_102_5_W0_en;
  wire  mem_102_5_W0_mask;
  wire [25:0] mem_102_6_R0_addr;
  wire  mem_102_6_R0_clk;
  wire [7:0] mem_102_6_R0_data;
  wire  mem_102_6_R0_en;
  wire [25:0] mem_102_6_W0_addr;
  wire  mem_102_6_W0_clk;
  wire [7:0] mem_102_6_W0_data;
  wire  mem_102_6_W0_en;
  wire  mem_102_6_W0_mask;
  wire [25:0] mem_102_7_R0_addr;
  wire  mem_102_7_R0_clk;
  wire [7:0] mem_102_7_R0_data;
  wire  mem_102_7_R0_en;
  wire [25:0] mem_102_7_W0_addr;
  wire  mem_102_7_W0_clk;
  wire [7:0] mem_102_7_W0_data;
  wire  mem_102_7_W0_en;
  wire  mem_102_7_W0_mask;
  wire [25:0] mem_103_0_R0_addr;
  wire  mem_103_0_R0_clk;
  wire [7:0] mem_103_0_R0_data;
  wire  mem_103_0_R0_en;
  wire [25:0] mem_103_0_W0_addr;
  wire  mem_103_0_W0_clk;
  wire [7:0] mem_103_0_W0_data;
  wire  mem_103_0_W0_en;
  wire  mem_103_0_W0_mask;
  wire [25:0] mem_103_1_R0_addr;
  wire  mem_103_1_R0_clk;
  wire [7:0] mem_103_1_R0_data;
  wire  mem_103_1_R0_en;
  wire [25:0] mem_103_1_W0_addr;
  wire  mem_103_1_W0_clk;
  wire [7:0] mem_103_1_W0_data;
  wire  mem_103_1_W0_en;
  wire  mem_103_1_W0_mask;
  wire [25:0] mem_103_2_R0_addr;
  wire  mem_103_2_R0_clk;
  wire [7:0] mem_103_2_R0_data;
  wire  mem_103_2_R0_en;
  wire [25:0] mem_103_2_W0_addr;
  wire  mem_103_2_W0_clk;
  wire [7:0] mem_103_2_W0_data;
  wire  mem_103_2_W0_en;
  wire  mem_103_2_W0_mask;
  wire [25:0] mem_103_3_R0_addr;
  wire  mem_103_3_R0_clk;
  wire [7:0] mem_103_3_R0_data;
  wire  mem_103_3_R0_en;
  wire [25:0] mem_103_3_W0_addr;
  wire  mem_103_3_W0_clk;
  wire [7:0] mem_103_3_W0_data;
  wire  mem_103_3_W0_en;
  wire  mem_103_3_W0_mask;
  wire [25:0] mem_103_4_R0_addr;
  wire  mem_103_4_R0_clk;
  wire [7:0] mem_103_4_R0_data;
  wire  mem_103_4_R0_en;
  wire [25:0] mem_103_4_W0_addr;
  wire  mem_103_4_W0_clk;
  wire [7:0] mem_103_4_W0_data;
  wire  mem_103_4_W0_en;
  wire  mem_103_4_W0_mask;
  wire [25:0] mem_103_5_R0_addr;
  wire  mem_103_5_R0_clk;
  wire [7:0] mem_103_5_R0_data;
  wire  mem_103_5_R0_en;
  wire [25:0] mem_103_5_W0_addr;
  wire  mem_103_5_W0_clk;
  wire [7:0] mem_103_5_W0_data;
  wire  mem_103_5_W0_en;
  wire  mem_103_5_W0_mask;
  wire [25:0] mem_103_6_R0_addr;
  wire  mem_103_6_R0_clk;
  wire [7:0] mem_103_6_R0_data;
  wire  mem_103_6_R0_en;
  wire [25:0] mem_103_6_W0_addr;
  wire  mem_103_6_W0_clk;
  wire [7:0] mem_103_6_W0_data;
  wire  mem_103_6_W0_en;
  wire  mem_103_6_W0_mask;
  wire [25:0] mem_103_7_R0_addr;
  wire  mem_103_7_R0_clk;
  wire [7:0] mem_103_7_R0_data;
  wire  mem_103_7_R0_en;
  wire [25:0] mem_103_7_W0_addr;
  wire  mem_103_7_W0_clk;
  wire [7:0] mem_103_7_W0_data;
  wire  mem_103_7_W0_en;
  wire  mem_103_7_W0_mask;
  wire [25:0] mem_104_0_R0_addr;
  wire  mem_104_0_R0_clk;
  wire [7:0] mem_104_0_R0_data;
  wire  mem_104_0_R0_en;
  wire [25:0] mem_104_0_W0_addr;
  wire  mem_104_0_W0_clk;
  wire [7:0] mem_104_0_W0_data;
  wire  mem_104_0_W0_en;
  wire  mem_104_0_W0_mask;
  wire [25:0] mem_104_1_R0_addr;
  wire  mem_104_1_R0_clk;
  wire [7:0] mem_104_1_R0_data;
  wire  mem_104_1_R0_en;
  wire [25:0] mem_104_1_W0_addr;
  wire  mem_104_1_W0_clk;
  wire [7:0] mem_104_1_W0_data;
  wire  mem_104_1_W0_en;
  wire  mem_104_1_W0_mask;
  wire [25:0] mem_104_2_R0_addr;
  wire  mem_104_2_R0_clk;
  wire [7:0] mem_104_2_R0_data;
  wire  mem_104_2_R0_en;
  wire [25:0] mem_104_2_W0_addr;
  wire  mem_104_2_W0_clk;
  wire [7:0] mem_104_2_W0_data;
  wire  mem_104_2_W0_en;
  wire  mem_104_2_W0_mask;
  wire [25:0] mem_104_3_R0_addr;
  wire  mem_104_3_R0_clk;
  wire [7:0] mem_104_3_R0_data;
  wire  mem_104_3_R0_en;
  wire [25:0] mem_104_3_W0_addr;
  wire  mem_104_3_W0_clk;
  wire [7:0] mem_104_3_W0_data;
  wire  mem_104_3_W0_en;
  wire  mem_104_3_W0_mask;
  wire [25:0] mem_104_4_R0_addr;
  wire  mem_104_4_R0_clk;
  wire [7:0] mem_104_4_R0_data;
  wire  mem_104_4_R0_en;
  wire [25:0] mem_104_4_W0_addr;
  wire  mem_104_4_W0_clk;
  wire [7:0] mem_104_4_W0_data;
  wire  mem_104_4_W0_en;
  wire  mem_104_4_W0_mask;
  wire [25:0] mem_104_5_R0_addr;
  wire  mem_104_5_R0_clk;
  wire [7:0] mem_104_5_R0_data;
  wire  mem_104_5_R0_en;
  wire [25:0] mem_104_5_W0_addr;
  wire  mem_104_5_W0_clk;
  wire [7:0] mem_104_5_W0_data;
  wire  mem_104_5_W0_en;
  wire  mem_104_5_W0_mask;
  wire [25:0] mem_104_6_R0_addr;
  wire  mem_104_6_R0_clk;
  wire [7:0] mem_104_6_R0_data;
  wire  mem_104_6_R0_en;
  wire [25:0] mem_104_6_W0_addr;
  wire  mem_104_6_W0_clk;
  wire [7:0] mem_104_6_W0_data;
  wire  mem_104_6_W0_en;
  wire  mem_104_6_W0_mask;
  wire [25:0] mem_104_7_R0_addr;
  wire  mem_104_7_R0_clk;
  wire [7:0] mem_104_7_R0_data;
  wire  mem_104_7_R0_en;
  wire [25:0] mem_104_7_W0_addr;
  wire  mem_104_7_W0_clk;
  wire [7:0] mem_104_7_W0_data;
  wire  mem_104_7_W0_en;
  wire  mem_104_7_W0_mask;
  wire [25:0] mem_105_0_R0_addr;
  wire  mem_105_0_R0_clk;
  wire [7:0] mem_105_0_R0_data;
  wire  mem_105_0_R0_en;
  wire [25:0] mem_105_0_W0_addr;
  wire  mem_105_0_W0_clk;
  wire [7:0] mem_105_0_W0_data;
  wire  mem_105_0_W0_en;
  wire  mem_105_0_W0_mask;
  wire [25:0] mem_105_1_R0_addr;
  wire  mem_105_1_R0_clk;
  wire [7:0] mem_105_1_R0_data;
  wire  mem_105_1_R0_en;
  wire [25:0] mem_105_1_W0_addr;
  wire  mem_105_1_W0_clk;
  wire [7:0] mem_105_1_W0_data;
  wire  mem_105_1_W0_en;
  wire  mem_105_1_W0_mask;
  wire [25:0] mem_105_2_R0_addr;
  wire  mem_105_2_R0_clk;
  wire [7:0] mem_105_2_R0_data;
  wire  mem_105_2_R0_en;
  wire [25:0] mem_105_2_W0_addr;
  wire  mem_105_2_W0_clk;
  wire [7:0] mem_105_2_W0_data;
  wire  mem_105_2_W0_en;
  wire  mem_105_2_W0_mask;
  wire [25:0] mem_105_3_R0_addr;
  wire  mem_105_3_R0_clk;
  wire [7:0] mem_105_3_R0_data;
  wire  mem_105_3_R0_en;
  wire [25:0] mem_105_3_W0_addr;
  wire  mem_105_3_W0_clk;
  wire [7:0] mem_105_3_W0_data;
  wire  mem_105_3_W0_en;
  wire  mem_105_3_W0_mask;
  wire [25:0] mem_105_4_R0_addr;
  wire  mem_105_4_R0_clk;
  wire [7:0] mem_105_4_R0_data;
  wire  mem_105_4_R0_en;
  wire [25:0] mem_105_4_W0_addr;
  wire  mem_105_4_W0_clk;
  wire [7:0] mem_105_4_W0_data;
  wire  mem_105_4_W0_en;
  wire  mem_105_4_W0_mask;
  wire [25:0] mem_105_5_R0_addr;
  wire  mem_105_5_R0_clk;
  wire [7:0] mem_105_5_R0_data;
  wire  mem_105_5_R0_en;
  wire [25:0] mem_105_5_W0_addr;
  wire  mem_105_5_W0_clk;
  wire [7:0] mem_105_5_W0_data;
  wire  mem_105_5_W0_en;
  wire  mem_105_5_W0_mask;
  wire [25:0] mem_105_6_R0_addr;
  wire  mem_105_6_R0_clk;
  wire [7:0] mem_105_6_R0_data;
  wire  mem_105_6_R0_en;
  wire [25:0] mem_105_6_W0_addr;
  wire  mem_105_6_W0_clk;
  wire [7:0] mem_105_6_W0_data;
  wire  mem_105_6_W0_en;
  wire  mem_105_6_W0_mask;
  wire [25:0] mem_105_7_R0_addr;
  wire  mem_105_7_R0_clk;
  wire [7:0] mem_105_7_R0_data;
  wire  mem_105_7_R0_en;
  wire [25:0] mem_105_7_W0_addr;
  wire  mem_105_7_W0_clk;
  wire [7:0] mem_105_7_W0_data;
  wire  mem_105_7_W0_en;
  wire  mem_105_7_W0_mask;
  wire [25:0] mem_106_0_R0_addr;
  wire  mem_106_0_R0_clk;
  wire [7:0] mem_106_0_R0_data;
  wire  mem_106_0_R0_en;
  wire [25:0] mem_106_0_W0_addr;
  wire  mem_106_0_W0_clk;
  wire [7:0] mem_106_0_W0_data;
  wire  mem_106_0_W0_en;
  wire  mem_106_0_W0_mask;
  wire [25:0] mem_106_1_R0_addr;
  wire  mem_106_1_R0_clk;
  wire [7:0] mem_106_1_R0_data;
  wire  mem_106_1_R0_en;
  wire [25:0] mem_106_1_W0_addr;
  wire  mem_106_1_W0_clk;
  wire [7:0] mem_106_1_W0_data;
  wire  mem_106_1_W0_en;
  wire  mem_106_1_W0_mask;
  wire [25:0] mem_106_2_R0_addr;
  wire  mem_106_2_R0_clk;
  wire [7:0] mem_106_2_R0_data;
  wire  mem_106_2_R0_en;
  wire [25:0] mem_106_2_W0_addr;
  wire  mem_106_2_W0_clk;
  wire [7:0] mem_106_2_W0_data;
  wire  mem_106_2_W0_en;
  wire  mem_106_2_W0_mask;
  wire [25:0] mem_106_3_R0_addr;
  wire  mem_106_3_R0_clk;
  wire [7:0] mem_106_3_R0_data;
  wire  mem_106_3_R0_en;
  wire [25:0] mem_106_3_W0_addr;
  wire  mem_106_3_W0_clk;
  wire [7:0] mem_106_3_W0_data;
  wire  mem_106_3_W0_en;
  wire  mem_106_3_W0_mask;
  wire [25:0] mem_106_4_R0_addr;
  wire  mem_106_4_R0_clk;
  wire [7:0] mem_106_4_R0_data;
  wire  mem_106_4_R0_en;
  wire [25:0] mem_106_4_W0_addr;
  wire  mem_106_4_W0_clk;
  wire [7:0] mem_106_4_W0_data;
  wire  mem_106_4_W0_en;
  wire  mem_106_4_W0_mask;
  wire [25:0] mem_106_5_R0_addr;
  wire  mem_106_5_R0_clk;
  wire [7:0] mem_106_5_R0_data;
  wire  mem_106_5_R0_en;
  wire [25:0] mem_106_5_W0_addr;
  wire  mem_106_5_W0_clk;
  wire [7:0] mem_106_5_W0_data;
  wire  mem_106_5_W0_en;
  wire  mem_106_5_W0_mask;
  wire [25:0] mem_106_6_R0_addr;
  wire  mem_106_6_R0_clk;
  wire [7:0] mem_106_6_R0_data;
  wire  mem_106_6_R0_en;
  wire [25:0] mem_106_6_W0_addr;
  wire  mem_106_6_W0_clk;
  wire [7:0] mem_106_6_W0_data;
  wire  mem_106_6_W0_en;
  wire  mem_106_6_W0_mask;
  wire [25:0] mem_106_7_R0_addr;
  wire  mem_106_7_R0_clk;
  wire [7:0] mem_106_7_R0_data;
  wire  mem_106_7_R0_en;
  wire [25:0] mem_106_7_W0_addr;
  wire  mem_106_7_W0_clk;
  wire [7:0] mem_106_7_W0_data;
  wire  mem_106_7_W0_en;
  wire  mem_106_7_W0_mask;
  wire [25:0] mem_107_0_R0_addr;
  wire  mem_107_0_R0_clk;
  wire [7:0] mem_107_0_R0_data;
  wire  mem_107_0_R0_en;
  wire [25:0] mem_107_0_W0_addr;
  wire  mem_107_0_W0_clk;
  wire [7:0] mem_107_0_W0_data;
  wire  mem_107_0_W0_en;
  wire  mem_107_0_W0_mask;
  wire [25:0] mem_107_1_R0_addr;
  wire  mem_107_1_R0_clk;
  wire [7:0] mem_107_1_R0_data;
  wire  mem_107_1_R0_en;
  wire [25:0] mem_107_1_W0_addr;
  wire  mem_107_1_W0_clk;
  wire [7:0] mem_107_1_W0_data;
  wire  mem_107_1_W0_en;
  wire  mem_107_1_W0_mask;
  wire [25:0] mem_107_2_R0_addr;
  wire  mem_107_2_R0_clk;
  wire [7:0] mem_107_2_R0_data;
  wire  mem_107_2_R0_en;
  wire [25:0] mem_107_2_W0_addr;
  wire  mem_107_2_W0_clk;
  wire [7:0] mem_107_2_W0_data;
  wire  mem_107_2_W0_en;
  wire  mem_107_2_W0_mask;
  wire [25:0] mem_107_3_R0_addr;
  wire  mem_107_3_R0_clk;
  wire [7:0] mem_107_3_R0_data;
  wire  mem_107_3_R0_en;
  wire [25:0] mem_107_3_W0_addr;
  wire  mem_107_3_W0_clk;
  wire [7:0] mem_107_3_W0_data;
  wire  mem_107_3_W0_en;
  wire  mem_107_3_W0_mask;
  wire [25:0] mem_107_4_R0_addr;
  wire  mem_107_4_R0_clk;
  wire [7:0] mem_107_4_R0_data;
  wire  mem_107_4_R0_en;
  wire [25:0] mem_107_4_W0_addr;
  wire  mem_107_4_W0_clk;
  wire [7:0] mem_107_4_W0_data;
  wire  mem_107_4_W0_en;
  wire  mem_107_4_W0_mask;
  wire [25:0] mem_107_5_R0_addr;
  wire  mem_107_5_R0_clk;
  wire [7:0] mem_107_5_R0_data;
  wire  mem_107_5_R0_en;
  wire [25:0] mem_107_5_W0_addr;
  wire  mem_107_5_W0_clk;
  wire [7:0] mem_107_5_W0_data;
  wire  mem_107_5_W0_en;
  wire  mem_107_5_W0_mask;
  wire [25:0] mem_107_6_R0_addr;
  wire  mem_107_6_R0_clk;
  wire [7:0] mem_107_6_R0_data;
  wire  mem_107_6_R0_en;
  wire [25:0] mem_107_6_W0_addr;
  wire  mem_107_6_W0_clk;
  wire [7:0] mem_107_6_W0_data;
  wire  mem_107_6_W0_en;
  wire  mem_107_6_W0_mask;
  wire [25:0] mem_107_7_R0_addr;
  wire  mem_107_7_R0_clk;
  wire [7:0] mem_107_7_R0_data;
  wire  mem_107_7_R0_en;
  wire [25:0] mem_107_7_W0_addr;
  wire  mem_107_7_W0_clk;
  wire [7:0] mem_107_7_W0_data;
  wire  mem_107_7_W0_en;
  wire  mem_107_7_W0_mask;
  wire [25:0] mem_108_0_R0_addr;
  wire  mem_108_0_R0_clk;
  wire [7:0] mem_108_0_R0_data;
  wire  mem_108_0_R0_en;
  wire [25:0] mem_108_0_W0_addr;
  wire  mem_108_0_W0_clk;
  wire [7:0] mem_108_0_W0_data;
  wire  mem_108_0_W0_en;
  wire  mem_108_0_W0_mask;
  wire [25:0] mem_108_1_R0_addr;
  wire  mem_108_1_R0_clk;
  wire [7:0] mem_108_1_R0_data;
  wire  mem_108_1_R0_en;
  wire [25:0] mem_108_1_W0_addr;
  wire  mem_108_1_W0_clk;
  wire [7:0] mem_108_1_W0_data;
  wire  mem_108_1_W0_en;
  wire  mem_108_1_W0_mask;
  wire [25:0] mem_108_2_R0_addr;
  wire  mem_108_2_R0_clk;
  wire [7:0] mem_108_2_R0_data;
  wire  mem_108_2_R0_en;
  wire [25:0] mem_108_2_W0_addr;
  wire  mem_108_2_W0_clk;
  wire [7:0] mem_108_2_W0_data;
  wire  mem_108_2_W0_en;
  wire  mem_108_2_W0_mask;
  wire [25:0] mem_108_3_R0_addr;
  wire  mem_108_3_R0_clk;
  wire [7:0] mem_108_3_R0_data;
  wire  mem_108_3_R0_en;
  wire [25:0] mem_108_3_W0_addr;
  wire  mem_108_3_W0_clk;
  wire [7:0] mem_108_3_W0_data;
  wire  mem_108_3_W0_en;
  wire  mem_108_3_W0_mask;
  wire [25:0] mem_108_4_R0_addr;
  wire  mem_108_4_R0_clk;
  wire [7:0] mem_108_4_R0_data;
  wire  mem_108_4_R0_en;
  wire [25:0] mem_108_4_W0_addr;
  wire  mem_108_4_W0_clk;
  wire [7:0] mem_108_4_W0_data;
  wire  mem_108_4_W0_en;
  wire  mem_108_4_W0_mask;
  wire [25:0] mem_108_5_R0_addr;
  wire  mem_108_5_R0_clk;
  wire [7:0] mem_108_5_R0_data;
  wire  mem_108_5_R0_en;
  wire [25:0] mem_108_5_W0_addr;
  wire  mem_108_5_W0_clk;
  wire [7:0] mem_108_5_W0_data;
  wire  mem_108_5_W0_en;
  wire  mem_108_5_W0_mask;
  wire [25:0] mem_108_6_R0_addr;
  wire  mem_108_6_R0_clk;
  wire [7:0] mem_108_6_R0_data;
  wire  mem_108_6_R0_en;
  wire [25:0] mem_108_6_W0_addr;
  wire  mem_108_6_W0_clk;
  wire [7:0] mem_108_6_W0_data;
  wire  mem_108_6_W0_en;
  wire  mem_108_6_W0_mask;
  wire [25:0] mem_108_7_R0_addr;
  wire  mem_108_7_R0_clk;
  wire [7:0] mem_108_7_R0_data;
  wire  mem_108_7_R0_en;
  wire [25:0] mem_108_7_W0_addr;
  wire  mem_108_7_W0_clk;
  wire [7:0] mem_108_7_W0_data;
  wire  mem_108_7_W0_en;
  wire  mem_108_7_W0_mask;
  wire [25:0] mem_109_0_R0_addr;
  wire  mem_109_0_R0_clk;
  wire [7:0] mem_109_0_R0_data;
  wire  mem_109_0_R0_en;
  wire [25:0] mem_109_0_W0_addr;
  wire  mem_109_0_W0_clk;
  wire [7:0] mem_109_0_W0_data;
  wire  mem_109_0_W0_en;
  wire  mem_109_0_W0_mask;
  wire [25:0] mem_109_1_R0_addr;
  wire  mem_109_1_R0_clk;
  wire [7:0] mem_109_1_R0_data;
  wire  mem_109_1_R0_en;
  wire [25:0] mem_109_1_W0_addr;
  wire  mem_109_1_W0_clk;
  wire [7:0] mem_109_1_W0_data;
  wire  mem_109_1_W0_en;
  wire  mem_109_1_W0_mask;
  wire [25:0] mem_109_2_R0_addr;
  wire  mem_109_2_R0_clk;
  wire [7:0] mem_109_2_R0_data;
  wire  mem_109_2_R0_en;
  wire [25:0] mem_109_2_W0_addr;
  wire  mem_109_2_W0_clk;
  wire [7:0] mem_109_2_W0_data;
  wire  mem_109_2_W0_en;
  wire  mem_109_2_W0_mask;
  wire [25:0] mem_109_3_R0_addr;
  wire  mem_109_3_R0_clk;
  wire [7:0] mem_109_3_R0_data;
  wire  mem_109_3_R0_en;
  wire [25:0] mem_109_3_W0_addr;
  wire  mem_109_3_W0_clk;
  wire [7:0] mem_109_3_W0_data;
  wire  mem_109_3_W0_en;
  wire  mem_109_3_W0_mask;
  wire [25:0] mem_109_4_R0_addr;
  wire  mem_109_4_R0_clk;
  wire [7:0] mem_109_4_R0_data;
  wire  mem_109_4_R0_en;
  wire [25:0] mem_109_4_W0_addr;
  wire  mem_109_4_W0_clk;
  wire [7:0] mem_109_4_W0_data;
  wire  mem_109_4_W0_en;
  wire  mem_109_4_W0_mask;
  wire [25:0] mem_109_5_R0_addr;
  wire  mem_109_5_R0_clk;
  wire [7:0] mem_109_5_R0_data;
  wire  mem_109_5_R0_en;
  wire [25:0] mem_109_5_W0_addr;
  wire  mem_109_5_W0_clk;
  wire [7:0] mem_109_5_W0_data;
  wire  mem_109_5_W0_en;
  wire  mem_109_5_W0_mask;
  wire [25:0] mem_109_6_R0_addr;
  wire  mem_109_6_R0_clk;
  wire [7:0] mem_109_6_R0_data;
  wire  mem_109_6_R0_en;
  wire [25:0] mem_109_6_W0_addr;
  wire  mem_109_6_W0_clk;
  wire [7:0] mem_109_6_W0_data;
  wire  mem_109_6_W0_en;
  wire  mem_109_6_W0_mask;
  wire [25:0] mem_109_7_R0_addr;
  wire  mem_109_7_R0_clk;
  wire [7:0] mem_109_7_R0_data;
  wire  mem_109_7_R0_en;
  wire [25:0] mem_109_7_W0_addr;
  wire  mem_109_7_W0_clk;
  wire [7:0] mem_109_7_W0_data;
  wire  mem_109_7_W0_en;
  wire  mem_109_7_W0_mask;
  wire [25:0] mem_110_0_R0_addr;
  wire  mem_110_0_R0_clk;
  wire [7:0] mem_110_0_R0_data;
  wire  mem_110_0_R0_en;
  wire [25:0] mem_110_0_W0_addr;
  wire  mem_110_0_W0_clk;
  wire [7:0] mem_110_0_W0_data;
  wire  mem_110_0_W0_en;
  wire  mem_110_0_W0_mask;
  wire [25:0] mem_110_1_R0_addr;
  wire  mem_110_1_R0_clk;
  wire [7:0] mem_110_1_R0_data;
  wire  mem_110_1_R0_en;
  wire [25:0] mem_110_1_W0_addr;
  wire  mem_110_1_W0_clk;
  wire [7:0] mem_110_1_W0_data;
  wire  mem_110_1_W0_en;
  wire  mem_110_1_W0_mask;
  wire [25:0] mem_110_2_R0_addr;
  wire  mem_110_2_R0_clk;
  wire [7:0] mem_110_2_R0_data;
  wire  mem_110_2_R0_en;
  wire [25:0] mem_110_2_W0_addr;
  wire  mem_110_2_W0_clk;
  wire [7:0] mem_110_2_W0_data;
  wire  mem_110_2_W0_en;
  wire  mem_110_2_W0_mask;
  wire [25:0] mem_110_3_R0_addr;
  wire  mem_110_3_R0_clk;
  wire [7:0] mem_110_3_R0_data;
  wire  mem_110_3_R0_en;
  wire [25:0] mem_110_3_W0_addr;
  wire  mem_110_3_W0_clk;
  wire [7:0] mem_110_3_W0_data;
  wire  mem_110_3_W0_en;
  wire  mem_110_3_W0_mask;
  wire [25:0] mem_110_4_R0_addr;
  wire  mem_110_4_R0_clk;
  wire [7:0] mem_110_4_R0_data;
  wire  mem_110_4_R0_en;
  wire [25:0] mem_110_4_W0_addr;
  wire  mem_110_4_W0_clk;
  wire [7:0] mem_110_4_W0_data;
  wire  mem_110_4_W0_en;
  wire  mem_110_4_W0_mask;
  wire [25:0] mem_110_5_R0_addr;
  wire  mem_110_5_R0_clk;
  wire [7:0] mem_110_5_R0_data;
  wire  mem_110_5_R0_en;
  wire [25:0] mem_110_5_W0_addr;
  wire  mem_110_5_W0_clk;
  wire [7:0] mem_110_5_W0_data;
  wire  mem_110_5_W0_en;
  wire  mem_110_5_W0_mask;
  wire [25:0] mem_110_6_R0_addr;
  wire  mem_110_6_R0_clk;
  wire [7:0] mem_110_6_R0_data;
  wire  mem_110_6_R0_en;
  wire [25:0] mem_110_6_W0_addr;
  wire  mem_110_6_W0_clk;
  wire [7:0] mem_110_6_W0_data;
  wire  mem_110_6_W0_en;
  wire  mem_110_6_W0_mask;
  wire [25:0] mem_110_7_R0_addr;
  wire  mem_110_7_R0_clk;
  wire [7:0] mem_110_7_R0_data;
  wire  mem_110_7_R0_en;
  wire [25:0] mem_110_7_W0_addr;
  wire  mem_110_7_W0_clk;
  wire [7:0] mem_110_7_W0_data;
  wire  mem_110_7_W0_en;
  wire  mem_110_7_W0_mask;
  wire [25:0] mem_111_0_R0_addr;
  wire  mem_111_0_R0_clk;
  wire [7:0] mem_111_0_R0_data;
  wire  mem_111_0_R0_en;
  wire [25:0] mem_111_0_W0_addr;
  wire  mem_111_0_W0_clk;
  wire [7:0] mem_111_0_W0_data;
  wire  mem_111_0_W0_en;
  wire  mem_111_0_W0_mask;
  wire [25:0] mem_111_1_R0_addr;
  wire  mem_111_1_R0_clk;
  wire [7:0] mem_111_1_R0_data;
  wire  mem_111_1_R0_en;
  wire [25:0] mem_111_1_W0_addr;
  wire  mem_111_1_W0_clk;
  wire [7:0] mem_111_1_W0_data;
  wire  mem_111_1_W0_en;
  wire  mem_111_1_W0_mask;
  wire [25:0] mem_111_2_R0_addr;
  wire  mem_111_2_R0_clk;
  wire [7:0] mem_111_2_R0_data;
  wire  mem_111_2_R0_en;
  wire [25:0] mem_111_2_W0_addr;
  wire  mem_111_2_W0_clk;
  wire [7:0] mem_111_2_W0_data;
  wire  mem_111_2_W0_en;
  wire  mem_111_2_W0_mask;
  wire [25:0] mem_111_3_R0_addr;
  wire  mem_111_3_R0_clk;
  wire [7:0] mem_111_3_R0_data;
  wire  mem_111_3_R0_en;
  wire [25:0] mem_111_3_W0_addr;
  wire  mem_111_3_W0_clk;
  wire [7:0] mem_111_3_W0_data;
  wire  mem_111_3_W0_en;
  wire  mem_111_3_W0_mask;
  wire [25:0] mem_111_4_R0_addr;
  wire  mem_111_4_R0_clk;
  wire [7:0] mem_111_4_R0_data;
  wire  mem_111_4_R0_en;
  wire [25:0] mem_111_4_W0_addr;
  wire  mem_111_4_W0_clk;
  wire [7:0] mem_111_4_W0_data;
  wire  mem_111_4_W0_en;
  wire  mem_111_4_W0_mask;
  wire [25:0] mem_111_5_R0_addr;
  wire  mem_111_5_R0_clk;
  wire [7:0] mem_111_5_R0_data;
  wire  mem_111_5_R0_en;
  wire [25:0] mem_111_5_W0_addr;
  wire  mem_111_5_W0_clk;
  wire [7:0] mem_111_5_W0_data;
  wire  mem_111_5_W0_en;
  wire  mem_111_5_W0_mask;
  wire [25:0] mem_111_6_R0_addr;
  wire  mem_111_6_R0_clk;
  wire [7:0] mem_111_6_R0_data;
  wire  mem_111_6_R0_en;
  wire [25:0] mem_111_6_W0_addr;
  wire  mem_111_6_W0_clk;
  wire [7:0] mem_111_6_W0_data;
  wire  mem_111_6_W0_en;
  wire  mem_111_6_W0_mask;
  wire [25:0] mem_111_7_R0_addr;
  wire  mem_111_7_R0_clk;
  wire [7:0] mem_111_7_R0_data;
  wire  mem_111_7_R0_en;
  wire [25:0] mem_111_7_W0_addr;
  wire  mem_111_7_W0_clk;
  wire [7:0] mem_111_7_W0_data;
  wire  mem_111_7_W0_en;
  wire  mem_111_7_W0_mask;
  wire [25:0] mem_112_0_R0_addr;
  wire  mem_112_0_R0_clk;
  wire [7:0] mem_112_0_R0_data;
  wire  mem_112_0_R0_en;
  wire [25:0] mem_112_0_W0_addr;
  wire  mem_112_0_W0_clk;
  wire [7:0] mem_112_0_W0_data;
  wire  mem_112_0_W0_en;
  wire  mem_112_0_W0_mask;
  wire [25:0] mem_112_1_R0_addr;
  wire  mem_112_1_R0_clk;
  wire [7:0] mem_112_1_R0_data;
  wire  mem_112_1_R0_en;
  wire [25:0] mem_112_1_W0_addr;
  wire  mem_112_1_W0_clk;
  wire [7:0] mem_112_1_W0_data;
  wire  mem_112_1_W0_en;
  wire  mem_112_1_W0_mask;
  wire [25:0] mem_112_2_R0_addr;
  wire  mem_112_2_R0_clk;
  wire [7:0] mem_112_2_R0_data;
  wire  mem_112_2_R0_en;
  wire [25:0] mem_112_2_W0_addr;
  wire  mem_112_2_W0_clk;
  wire [7:0] mem_112_2_W0_data;
  wire  mem_112_2_W0_en;
  wire  mem_112_2_W0_mask;
  wire [25:0] mem_112_3_R0_addr;
  wire  mem_112_3_R0_clk;
  wire [7:0] mem_112_3_R0_data;
  wire  mem_112_3_R0_en;
  wire [25:0] mem_112_3_W0_addr;
  wire  mem_112_3_W0_clk;
  wire [7:0] mem_112_3_W0_data;
  wire  mem_112_3_W0_en;
  wire  mem_112_3_W0_mask;
  wire [25:0] mem_112_4_R0_addr;
  wire  mem_112_4_R0_clk;
  wire [7:0] mem_112_4_R0_data;
  wire  mem_112_4_R0_en;
  wire [25:0] mem_112_4_W0_addr;
  wire  mem_112_4_W0_clk;
  wire [7:0] mem_112_4_W0_data;
  wire  mem_112_4_W0_en;
  wire  mem_112_4_W0_mask;
  wire [25:0] mem_112_5_R0_addr;
  wire  mem_112_5_R0_clk;
  wire [7:0] mem_112_5_R0_data;
  wire  mem_112_5_R0_en;
  wire [25:0] mem_112_5_W0_addr;
  wire  mem_112_5_W0_clk;
  wire [7:0] mem_112_5_W0_data;
  wire  mem_112_5_W0_en;
  wire  mem_112_5_W0_mask;
  wire [25:0] mem_112_6_R0_addr;
  wire  mem_112_6_R0_clk;
  wire [7:0] mem_112_6_R0_data;
  wire  mem_112_6_R0_en;
  wire [25:0] mem_112_6_W0_addr;
  wire  mem_112_6_W0_clk;
  wire [7:0] mem_112_6_W0_data;
  wire  mem_112_6_W0_en;
  wire  mem_112_6_W0_mask;
  wire [25:0] mem_112_7_R0_addr;
  wire  mem_112_7_R0_clk;
  wire [7:0] mem_112_7_R0_data;
  wire  mem_112_7_R0_en;
  wire [25:0] mem_112_7_W0_addr;
  wire  mem_112_7_W0_clk;
  wire [7:0] mem_112_7_W0_data;
  wire  mem_112_7_W0_en;
  wire  mem_112_7_W0_mask;
  wire [25:0] mem_113_0_R0_addr;
  wire  mem_113_0_R0_clk;
  wire [7:0] mem_113_0_R0_data;
  wire  mem_113_0_R0_en;
  wire [25:0] mem_113_0_W0_addr;
  wire  mem_113_0_W0_clk;
  wire [7:0] mem_113_0_W0_data;
  wire  mem_113_0_W0_en;
  wire  mem_113_0_W0_mask;
  wire [25:0] mem_113_1_R0_addr;
  wire  mem_113_1_R0_clk;
  wire [7:0] mem_113_1_R0_data;
  wire  mem_113_1_R0_en;
  wire [25:0] mem_113_1_W0_addr;
  wire  mem_113_1_W0_clk;
  wire [7:0] mem_113_1_W0_data;
  wire  mem_113_1_W0_en;
  wire  mem_113_1_W0_mask;
  wire [25:0] mem_113_2_R0_addr;
  wire  mem_113_2_R0_clk;
  wire [7:0] mem_113_2_R0_data;
  wire  mem_113_2_R0_en;
  wire [25:0] mem_113_2_W0_addr;
  wire  mem_113_2_W0_clk;
  wire [7:0] mem_113_2_W0_data;
  wire  mem_113_2_W0_en;
  wire  mem_113_2_W0_mask;
  wire [25:0] mem_113_3_R0_addr;
  wire  mem_113_3_R0_clk;
  wire [7:0] mem_113_3_R0_data;
  wire  mem_113_3_R0_en;
  wire [25:0] mem_113_3_W0_addr;
  wire  mem_113_3_W0_clk;
  wire [7:0] mem_113_3_W0_data;
  wire  mem_113_3_W0_en;
  wire  mem_113_3_W0_mask;
  wire [25:0] mem_113_4_R0_addr;
  wire  mem_113_4_R0_clk;
  wire [7:0] mem_113_4_R0_data;
  wire  mem_113_4_R0_en;
  wire [25:0] mem_113_4_W0_addr;
  wire  mem_113_4_W0_clk;
  wire [7:0] mem_113_4_W0_data;
  wire  mem_113_4_W0_en;
  wire  mem_113_4_W0_mask;
  wire [25:0] mem_113_5_R0_addr;
  wire  mem_113_5_R0_clk;
  wire [7:0] mem_113_5_R0_data;
  wire  mem_113_5_R0_en;
  wire [25:0] mem_113_5_W0_addr;
  wire  mem_113_5_W0_clk;
  wire [7:0] mem_113_5_W0_data;
  wire  mem_113_5_W0_en;
  wire  mem_113_5_W0_mask;
  wire [25:0] mem_113_6_R0_addr;
  wire  mem_113_6_R0_clk;
  wire [7:0] mem_113_6_R0_data;
  wire  mem_113_6_R0_en;
  wire [25:0] mem_113_6_W0_addr;
  wire  mem_113_6_W0_clk;
  wire [7:0] mem_113_6_W0_data;
  wire  mem_113_6_W0_en;
  wire  mem_113_6_W0_mask;
  wire [25:0] mem_113_7_R0_addr;
  wire  mem_113_7_R0_clk;
  wire [7:0] mem_113_7_R0_data;
  wire  mem_113_7_R0_en;
  wire [25:0] mem_113_7_W0_addr;
  wire  mem_113_7_W0_clk;
  wire [7:0] mem_113_7_W0_data;
  wire  mem_113_7_W0_en;
  wire  mem_113_7_W0_mask;
  wire [25:0] mem_114_0_R0_addr;
  wire  mem_114_0_R0_clk;
  wire [7:0] mem_114_0_R0_data;
  wire  mem_114_0_R0_en;
  wire [25:0] mem_114_0_W0_addr;
  wire  mem_114_0_W0_clk;
  wire [7:0] mem_114_0_W0_data;
  wire  mem_114_0_W0_en;
  wire  mem_114_0_W0_mask;
  wire [25:0] mem_114_1_R0_addr;
  wire  mem_114_1_R0_clk;
  wire [7:0] mem_114_1_R0_data;
  wire  mem_114_1_R0_en;
  wire [25:0] mem_114_1_W0_addr;
  wire  mem_114_1_W0_clk;
  wire [7:0] mem_114_1_W0_data;
  wire  mem_114_1_W0_en;
  wire  mem_114_1_W0_mask;
  wire [25:0] mem_114_2_R0_addr;
  wire  mem_114_2_R0_clk;
  wire [7:0] mem_114_2_R0_data;
  wire  mem_114_2_R0_en;
  wire [25:0] mem_114_2_W0_addr;
  wire  mem_114_2_W0_clk;
  wire [7:0] mem_114_2_W0_data;
  wire  mem_114_2_W0_en;
  wire  mem_114_2_W0_mask;
  wire [25:0] mem_114_3_R0_addr;
  wire  mem_114_3_R0_clk;
  wire [7:0] mem_114_3_R0_data;
  wire  mem_114_3_R0_en;
  wire [25:0] mem_114_3_W0_addr;
  wire  mem_114_3_W0_clk;
  wire [7:0] mem_114_3_W0_data;
  wire  mem_114_3_W0_en;
  wire  mem_114_3_W0_mask;
  wire [25:0] mem_114_4_R0_addr;
  wire  mem_114_4_R0_clk;
  wire [7:0] mem_114_4_R0_data;
  wire  mem_114_4_R0_en;
  wire [25:0] mem_114_4_W0_addr;
  wire  mem_114_4_W0_clk;
  wire [7:0] mem_114_4_W0_data;
  wire  mem_114_4_W0_en;
  wire  mem_114_4_W0_mask;
  wire [25:0] mem_114_5_R0_addr;
  wire  mem_114_5_R0_clk;
  wire [7:0] mem_114_5_R0_data;
  wire  mem_114_5_R0_en;
  wire [25:0] mem_114_5_W0_addr;
  wire  mem_114_5_W0_clk;
  wire [7:0] mem_114_5_W0_data;
  wire  mem_114_5_W0_en;
  wire  mem_114_5_W0_mask;
  wire [25:0] mem_114_6_R0_addr;
  wire  mem_114_6_R0_clk;
  wire [7:0] mem_114_6_R0_data;
  wire  mem_114_6_R0_en;
  wire [25:0] mem_114_6_W0_addr;
  wire  mem_114_6_W0_clk;
  wire [7:0] mem_114_6_W0_data;
  wire  mem_114_6_W0_en;
  wire  mem_114_6_W0_mask;
  wire [25:0] mem_114_7_R0_addr;
  wire  mem_114_7_R0_clk;
  wire [7:0] mem_114_7_R0_data;
  wire  mem_114_7_R0_en;
  wire [25:0] mem_114_7_W0_addr;
  wire  mem_114_7_W0_clk;
  wire [7:0] mem_114_7_W0_data;
  wire  mem_114_7_W0_en;
  wire  mem_114_7_W0_mask;
  wire [25:0] mem_115_0_R0_addr;
  wire  mem_115_0_R0_clk;
  wire [7:0] mem_115_0_R0_data;
  wire  mem_115_0_R0_en;
  wire [25:0] mem_115_0_W0_addr;
  wire  mem_115_0_W0_clk;
  wire [7:0] mem_115_0_W0_data;
  wire  mem_115_0_W0_en;
  wire  mem_115_0_W0_mask;
  wire [25:0] mem_115_1_R0_addr;
  wire  mem_115_1_R0_clk;
  wire [7:0] mem_115_1_R0_data;
  wire  mem_115_1_R0_en;
  wire [25:0] mem_115_1_W0_addr;
  wire  mem_115_1_W0_clk;
  wire [7:0] mem_115_1_W0_data;
  wire  mem_115_1_W0_en;
  wire  mem_115_1_W0_mask;
  wire [25:0] mem_115_2_R0_addr;
  wire  mem_115_2_R0_clk;
  wire [7:0] mem_115_2_R0_data;
  wire  mem_115_2_R0_en;
  wire [25:0] mem_115_2_W0_addr;
  wire  mem_115_2_W0_clk;
  wire [7:0] mem_115_2_W0_data;
  wire  mem_115_2_W0_en;
  wire  mem_115_2_W0_mask;
  wire [25:0] mem_115_3_R0_addr;
  wire  mem_115_3_R0_clk;
  wire [7:0] mem_115_3_R0_data;
  wire  mem_115_3_R0_en;
  wire [25:0] mem_115_3_W0_addr;
  wire  mem_115_3_W0_clk;
  wire [7:0] mem_115_3_W0_data;
  wire  mem_115_3_W0_en;
  wire  mem_115_3_W0_mask;
  wire [25:0] mem_115_4_R0_addr;
  wire  mem_115_4_R0_clk;
  wire [7:0] mem_115_4_R0_data;
  wire  mem_115_4_R0_en;
  wire [25:0] mem_115_4_W0_addr;
  wire  mem_115_4_W0_clk;
  wire [7:0] mem_115_4_W0_data;
  wire  mem_115_4_W0_en;
  wire  mem_115_4_W0_mask;
  wire [25:0] mem_115_5_R0_addr;
  wire  mem_115_5_R0_clk;
  wire [7:0] mem_115_5_R0_data;
  wire  mem_115_5_R0_en;
  wire [25:0] mem_115_5_W0_addr;
  wire  mem_115_5_W0_clk;
  wire [7:0] mem_115_5_W0_data;
  wire  mem_115_5_W0_en;
  wire  mem_115_5_W0_mask;
  wire [25:0] mem_115_6_R0_addr;
  wire  mem_115_6_R0_clk;
  wire [7:0] mem_115_6_R0_data;
  wire  mem_115_6_R0_en;
  wire [25:0] mem_115_6_W0_addr;
  wire  mem_115_6_W0_clk;
  wire [7:0] mem_115_6_W0_data;
  wire  mem_115_6_W0_en;
  wire  mem_115_6_W0_mask;
  wire [25:0] mem_115_7_R0_addr;
  wire  mem_115_7_R0_clk;
  wire [7:0] mem_115_7_R0_data;
  wire  mem_115_7_R0_en;
  wire [25:0] mem_115_7_W0_addr;
  wire  mem_115_7_W0_clk;
  wire [7:0] mem_115_7_W0_data;
  wire  mem_115_7_W0_en;
  wire  mem_115_7_W0_mask;
  wire [25:0] mem_116_0_R0_addr;
  wire  mem_116_0_R0_clk;
  wire [7:0] mem_116_0_R0_data;
  wire  mem_116_0_R0_en;
  wire [25:0] mem_116_0_W0_addr;
  wire  mem_116_0_W0_clk;
  wire [7:0] mem_116_0_W0_data;
  wire  mem_116_0_W0_en;
  wire  mem_116_0_W0_mask;
  wire [25:0] mem_116_1_R0_addr;
  wire  mem_116_1_R0_clk;
  wire [7:0] mem_116_1_R0_data;
  wire  mem_116_1_R0_en;
  wire [25:0] mem_116_1_W0_addr;
  wire  mem_116_1_W0_clk;
  wire [7:0] mem_116_1_W0_data;
  wire  mem_116_1_W0_en;
  wire  mem_116_1_W0_mask;
  wire [25:0] mem_116_2_R0_addr;
  wire  mem_116_2_R0_clk;
  wire [7:0] mem_116_2_R0_data;
  wire  mem_116_2_R0_en;
  wire [25:0] mem_116_2_W0_addr;
  wire  mem_116_2_W0_clk;
  wire [7:0] mem_116_2_W0_data;
  wire  mem_116_2_W0_en;
  wire  mem_116_2_W0_mask;
  wire [25:0] mem_116_3_R0_addr;
  wire  mem_116_3_R0_clk;
  wire [7:0] mem_116_3_R0_data;
  wire  mem_116_3_R0_en;
  wire [25:0] mem_116_3_W0_addr;
  wire  mem_116_3_W0_clk;
  wire [7:0] mem_116_3_W0_data;
  wire  mem_116_3_W0_en;
  wire  mem_116_3_W0_mask;
  wire [25:0] mem_116_4_R0_addr;
  wire  mem_116_4_R0_clk;
  wire [7:0] mem_116_4_R0_data;
  wire  mem_116_4_R0_en;
  wire [25:0] mem_116_4_W0_addr;
  wire  mem_116_4_W0_clk;
  wire [7:0] mem_116_4_W0_data;
  wire  mem_116_4_W0_en;
  wire  mem_116_4_W0_mask;
  wire [25:0] mem_116_5_R0_addr;
  wire  mem_116_5_R0_clk;
  wire [7:0] mem_116_5_R0_data;
  wire  mem_116_5_R0_en;
  wire [25:0] mem_116_5_W0_addr;
  wire  mem_116_5_W0_clk;
  wire [7:0] mem_116_5_W0_data;
  wire  mem_116_5_W0_en;
  wire  mem_116_5_W0_mask;
  wire [25:0] mem_116_6_R0_addr;
  wire  mem_116_6_R0_clk;
  wire [7:0] mem_116_6_R0_data;
  wire  mem_116_6_R0_en;
  wire [25:0] mem_116_6_W0_addr;
  wire  mem_116_6_W0_clk;
  wire [7:0] mem_116_6_W0_data;
  wire  mem_116_6_W0_en;
  wire  mem_116_6_W0_mask;
  wire [25:0] mem_116_7_R0_addr;
  wire  mem_116_7_R0_clk;
  wire [7:0] mem_116_7_R0_data;
  wire  mem_116_7_R0_en;
  wire [25:0] mem_116_7_W0_addr;
  wire  mem_116_7_W0_clk;
  wire [7:0] mem_116_7_W0_data;
  wire  mem_116_7_W0_en;
  wire  mem_116_7_W0_mask;
  wire [25:0] mem_117_0_R0_addr;
  wire  mem_117_0_R0_clk;
  wire [7:0] mem_117_0_R0_data;
  wire  mem_117_0_R0_en;
  wire [25:0] mem_117_0_W0_addr;
  wire  mem_117_0_W0_clk;
  wire [7:0] mem_117_0_W0_data;
  wire  mem_117_0_W0_en;
  wire  mem_117_0_W0_mask;
  wire [25:0] mem_117_1_R0_addr;
  wire  mem_117_1_R0_clk;
  wire [7:0] mem_117_1_R0_data;
  wire  mem_117_1_R0_en;
  wire [25:0] mem_117_1_W0_addr;
  wire  mem_117_1_W0_clk;
  wire [7:0] mem_117_1_W0_data;
  wire  mem_117_1_W0_en;
  wire  mem_117_1_W0_mask;
  wire [25:0] mem_117_2_R0_addr;
  wire  mem_117_2_R0_clk;
  wire [7:0] mem_117_2_R0_data;
  wire  mem_117_2_R0_en;
  wire [25:0] mem_117_2_W0_addr;
  wire  mem_117_2_W0_clk;
  wire [7:0] mem_117_2_W0_data;
  wire  mem_117_2_W0_en;
  wire  mem_117_2_W0_mask;
  wire [25:0] mem_117_3_R0_addr;
  wire  mem_117_3_R0_clk;
  wire [7:0] mem_117_3_R0_data;
  wire  mem_117_3_R0_en;
  wire [25:0] mem_117_3_W0_addr;
  wire  mem_117_3_W0_clk;
  wire [7:0] mem_117_3_W0_data;
  wire  mem_117_3_W0_en;
  wire  mem_117_3_W0_mask;
  wire [25:0] mem_117_4_R0_addr;
  wire  mem_117_4_R0_clk;
  wire [7:0] mem_117_4_R0_data;
  wire  mem_117_4_R0_en;
  wire [25:0] mem_117_4_W0_addr;
  wire  mem_117_4_W0_clk;
  wire [7:0] mem_117_4_W0_data;
  wire  mem_117_4_W0_en;
  wire  mem_117_4_W0_mask;
  wire [25:0] mem_117_5_R0_addr;
  wire  mem_117_5_R0_clk;
  wire [7:0] mem_117_5_R0_data;
  wire  mem_117_5_R0_en;
  wire [25:0] mem_117_5_W0_addr;
  wire  mem_117_5_W0_clk;
  wire [7:0] mem_117_5_W0_data;
  wire  mem_117_5_W0_en;
  wire  mem_117_5_W0_mask;
  wire [25:0] mem_117_6_R0_addr;
  wire  mem_117_6_R0_clk;
  wire [7:0] mem_117_6_R0_data;
  wire  mem_117_6_R0_en;
  wire [25:0] mem_117_6_W0_addr;
  wire  mem_117_6_W0_clk;
  wire [7:0] mem_117_6_W0_data;
  wire  mem_117_6_W0_en;
  wire  mem_117_6_W0_mask;
  wire [25:0] mem_117_7_R0_addr;
  wire  mem_117_7_R0_clk;
  wire [7:0] mem_117_7_R0_data;
  wire  mem_117_7_R0_en;
  wire [25:0] mem_117_7_W0_addr;
  wire  mem_117_7_W0_clk;
  wire [7:0] mem_117_7_W0_data;
  wire  mem_117_7_W0_en;
  wire  mem_117_7_W0_mask;
  wire [25:0] mem_118_0_R0_addr;
  wire  mem_118_0_R0_clk;
  wire [7:0] mem_118_0_R0_data;
  wire  mem_118_0_R0_en;
  wire [25:0] mem_118_0_W0_addr;
  wire  mem_118_0_W0_clk;
  wire [7:0] mem_118_0_W0_data;
  wire  mem_118_0_W0_en;
  wire  mem_118_0_W0_mask;
  wire [25:0] mem_118_1_R0_addr;
  wire  mem_118_1_R0_clk;
  wire [7:0] mem_118_1_R0_data;
  wire  mem_118_1_R0_en;
  wire [25:0] mem_118_1_W0_addr;
  wire  mem_118_1_W0_clk;
  wire [7:0] mem_118_1_W0_data;
  wire  mem_118_1_W0_en;
  wire  mem_118_1_W0_mask;
  wire [25:0] mem_118_2_R0_addr;
  wire  mem_118_2_R0_clk;
  wire [7:0] mem_118_2_R0_data;
  wire  mem_118_2_R0_en;
  wire [25:0] mem_118_2_W0_addr;
  wire  mem_118_2_W0_clk;
  wire [7:0] mem_118_2_W0_data;
  wire  mem_118_2_W0_en;
  wire  mem_118_2_W0_mask;
  wire [25:0] mem_118_3_R0_addr;
  wire  mem_118_3_R0_clk;
  wire [7:0] mem_118_3_R0_data;
  wire  mem_118_3_R0_en;
  wire [25:0] mem_118_3_W0_addr;
  wire  mem_118_3_W0_clk;
  wire [7:0] mem_118_3_W0_data;
  wire  mem_118_3_W0_en;
  wire  mem_118_3_W0_mask;
  wire [25:0] mem_118_4_R0_addr;
  wire  mem_118_4_R0_clk;
  wire [7:0] mem_118_4_R0_data;
  wire  mem_118_4_R0_en;
  wire [25:0] mem_118_4_W0_addr;
  wire  mem_118_4_W0_clk;
  wire [7:0] mem_118_4_W0_data;
  wire  mem_118_4_W0_en;
  wire  mem_118_4_W0_mask;
  wire [25:0] mem_118_5_R0_addr;
  wire  mem_118_5_R0_clk;
  wire [7:0] mem_118_5_R0_data;
  wire  mem_118_5_R0_en;
  wire [25:0] mem_118_5_W0_addr;
  wire  mem_118_5_W0_clk;
  wire [7:0] mem_118_5_W0_data;
  wire  mem_118_5_W0_en;
  wire  mem_118_5_W0_mask;
  wire [25:0] mem_118_6_R0_addr;
  wire  mem_118_6_R0_clk;
  wire [7:0] mem_118_6_R0_data;
  wire  mem_118_6_R0_en;
  wire [25:0] mem_118_6_W0_addr;
  wire  mem_118_6_W0_clk;
  wire [7:0] mem_118_6_W0_data;
  wire  mem_118_6_W0_en;
  wire  mem_118_6_W0_mask;
  wire [25:0] mem_118_7_R0_addr;
  wire  mem_118_7_R0_clk;
  wire [7:0] mem_118_7_R0_data;
  wire  mem_118_7_R0_en;
  wire [25:0] mem_118_7_W0_addr;
  wire  mem_118_7_W0_clk;
  wire [7:0] mem_118_7_W0_data;
  wire  mem_118_7_W0_en;
  wire  mem_118_7_W0_mask;
  wire [25:0] mem_119_0_R0_addr;
  wire  mem_119_0_R0_clk;
  wire [7:0] mem_119_0_R0_data;
  wire  mem_119_0_R0_en;
  wire [25:0] mem_119_0_W0_addr;
  wire  mem_119_0_W0_clk;
  wire [7:0] mem_119_0_W0_data;
  wire  mem_119_0_W0_en;
  wire  mem_119_0_W0_mask;
  wire [25:0] mem_119_1_R0_addr;
  wire  mem_119_1_R0_clk;
  wire [7:0] mem_119_1_R0_data;
  wire  mem_119_1_R0_en;
  wire [25:0] mem_119_1_W0_addr;
  wire  mem_119_1_W0_clk;
  wire [7:0] mem_119_1_W0_data;
  wire  mem_119_1_W0_en;
  wire  mem_119_1_W0_mask;
  wire [25:0] mem_119_2_R0_addr;
  wire  mem_119_2_R0_clk;
  wire [7:0] mem_119_2_R0_data;
  wire  mem_119_2_R0_en;
  wire [25:0] mem_119_2_W0_addr;
  wire  mem_119_2_W0_clk;
  wire [7:0] mem_119_2_W0_data;
  wire  mem_119_2_W0_en;
  wire  mem_119_2_W0_mask;
  wire [25:0] mem_119_3_R0_addr;
  wire  mem_119_3_R0_clk;
  wire [7:0] mem_119_3_R0_data;
  wire  mem_119_3_R0_en;
  wire [25:0] mem_119_3_W0_addr;
  wire  mem_119_3_W0_clk;
  wire [7:0] mem_119_3_W0_data;
  wire  mem_119_3_W0_en;
  wire  mem_119_3_W0_mask;
  wire [25:0] mem_119_4_R0_addr;
  wire  mem_119_4_R0_clk;
  wire [7:0] mem_119_4_R0_data;
  wire  mem_119_4_R0_en;
  wire [25:0] mem_119_4_W0_addr;
  wire  mem_119_4_W0_clk;
  wire [7:0] mem_119_4_W0_data;
  wire  mem_119_4_W0_en;
  wire  mem_119_4_W0_mask;
  wire [25:0] mem_119_5_R0_addr;
  wire  mem_119_5_R0_clk;
  wire [7:0] mem_119_5_R0_data;
  wire  mem_119_5_R0_en;
  wire [25:0] mem_119_5_W0_addr;
  wire  mem_119_5_W0_clk;
  wire [7:0] mem_119_5_W0_data;
  wire  mem_119_5_W0_en;
  wire  mem_119_5_W0_mask;
  wire [25:0] mem_119_6_R0_addr;
  wire  mem_119_6_R0_clk;
  wire [7:0] mem_119_6_R0_data;
  wire  mem_119_6_R0_en;
  wire [25:0] mem_119_6_W0_addr;
  wire  mem_119_6_W0_clk;
  wire [7:0] mem_119_6_W0_data;
  wire  mem_119_6_W0_en;
  wire  mem_119_6_W0_mask;
  wire [25:0] mem_119_7_R0_addr;
  wire  mem_119_7_R0_clk;
  wire [7:0] mem_119_7_R0_data;
  wire  mem_119_7_R0_en;
  wire [25:0] mem_119_7_W0_addr;
  wire  mem_119_7_W0_clk;
  wire [7:0] mem_119_7_W0_data;
  wire  mem_119_7_W0_en;
  wire  mem_119_7_W0_mask;
  wire [25:0] mem_120_0_R0_addr;
  wire  mem_120_0_R0_clk;
  wire [7:0] mem_120_0_R0_data;
  wire  mem_120_0_R0_en;
  wire [25:0] mem_120_0_W0_addr;
  wire  mem_120_0_W0_clk;
  wire [7:0] mem_120_0_W0_data;
  wire  mem_120_0_W0_en;
  wire  mem_120_0_W0_mask;
  wire [25:0] mem_120_1_R0_addr;
  wire  mem_120_1_R0_clk;
  wire [7:0] mem_120_1_R0_data;
  wire  mem_120_1_R0_en;
  wire [25:0] mem_120_1_W0_addr;
  wire  mem_120_1_W0_clk;
  wire [7:0] mem_120_1_W0_data;
  wire  mem_120_1_W0_en;
  wire  mem_120_1_W0_mask;
  wire [25:0] mem_120_2_R0_addr;
  wire  mem_120_2_R0_clk;
  wire [7:0] mem_120_2_R0_data;
  wire  mem_120_2_R0_en;
  wire [25:0] mem_120_2_W0_addr;
  wire  mem_120_2_W0_clk;
  wire [7:0] mem_120_2_W0_data;
  wire  mem_120_2_W0_en;
  wire  mem_120_2_W0_mask;
  wire [25:0] mem_120_3_R0_addr;
  wire  mem_120_3_R0_clk;
  wire [7:0] mem_120_3_R0_data;
  wire  mem_120_3_R0_en;
  wire [25:0] mem_120_3_W0_addr;
  wire  mem_120_3_W0_clk;
  wire [7:0] mem_120_3_W0_data;
  wire  mem_120_3_W0_en;
  wire  mem_120_3_W0_mask;
  wire [25:0] mem_120_4_R0_addr;
  wire  mem_120_4_R0_clk;
  wire [7:0] mem_120_4_R0_data;
  wire  mem_120_4_R0_en;
  wire [25:0] mem_120_4_W0_addr;
  wire  mem_120_4_W0_clk;
  wire [7:0] mem_120_4_W0_data;
  wire  mem_120_4_W0_en;
  wire  mem_120_4_W0_mask;
  wire [25:0] mem_120_5_R0_addr;
  wire  mem_120_5_R0_clk;
  wire [7:0] mem_120_5_R0_data;
  wire  mem_120_5_R0_en;
  wire [25:0] mem_120_5_W0_addr;
  wire  mem_120_5_W0_clk;
  wire [7:0] mem_120_5_W0_data;
  wire  mem_120_5_W0_en;
  wire  mem_120_5_W0_mask;
  wire [25:0] mem_120_6_R0_addr;
  wire  mem_120_6_R0_clk;
  wire [7:0] mem_120_6_R0_data;
  wire  mem_120_6_R0_en;
  wire [25:0] mem_120_6_W0_addr;
  wire  mem_120_6_W0_clk;
  wire [7:0] mem_120_6_W0_data;
  wire  mem_120_6_W0_en;
  wire  mem_120_6_W0_mask;
  wire [25:0] mem_120_7_R0_addr;
  wire  mem_120_7_R0_clk;
  wire [7:0] mem_120_7_R0_data;
  wire  mem_120_7_R0_en;
  wire [25:0] mem_120_7_W0_addr;
  wire  mem_120_7_W0_clk;
  wire [7:0] mem_120_7_W0_data;
  wire  mem_120_7_W0_en;
  wire  mem_120_7_W0_mask;
  wire [25:0] mem_121_0_R0_addr;
  wire  mem_121_0_R0_clk;
  wire [7:0] mem_121_0_R0_data;
  wire  mem_121_0_R0_en;
  wire [25:0] mem_121_0_W0_addr;
  wire  mem_121_0_W0_clk;
  wire [7:0] mem_121_0_W0_data;
  wire  mem_121_0_W0_en;
  wire  mem_121_0_W0_mask;
  wire [25:0] mem_121_1_R0_addr;
  wire  mem_121_1_R0_clk;
  wire [7:0] mem_121_1_R0_data;
  wire  mem_121_1_R0_en;
  wire [25:0] mem_121_1_W0_addr;
  wire  mem_121_1_W0_clk;
  wire [7:0] mem_121_1_W0_data;
  wire  mem_121_1_W0_en;
  wire  mem_121_1_W0_mask;
  wire [25:0] mem_121_2_R0_addr;
  wire  mem_121_2_R0_clk;
  wire [7:0] mem_121_2_R0_data;
  wire  mem_121_2_R0_en;
  wire [25:0] mem_121_2_W0_addr;
  wire  mem_121_2_W0_clk;
  wire [7:0] mem_121_2_W0_data;
  wire  mem_121_2_W0_en;
  wire  mem_121_2_W0_mask;
  wire [25:0] mem_121_3_R0_addr;
  wire  mem_121_3_R0_clk;
  wire [7:0] mem_121_3_R0_data;
  wire  mem_121_3_R0_en;
  wire [25:0] mem_121_3_W0_addr;
  wire  mem_121_3_W0_clk;
  wire [7:0] mem_121_3_W0_data;
  wire  mem_121_3_W0_en;
  wire  mem_121_3_W0_mask;
  wire [25:0] mem_121_4_R0_addr;
  wire  mem_121_4_R0_clk;
  wire [7:0] mem_121_4_R0_data;
  wire  mem_121_4_R0_en;
  wire [25:0] mem_121_4_W0_addr;
  wire  mem_121_4_W0_clk;
  wire [7:0] mem_121_4_W0_data;
  wire  mem_121_4_W0_en;
  wire  mem_121_4_W0_mask;
  wire [25:0] mem_121_5_R0_addr;
  wire  mem_121_5_R0_clk;
  wire [7:0] mem_121_5_R0_data;
  wire  mem_121_5_R0_en;
  wire [25:0] mem_121_5_W0_addr;
  wire  mem_121_5_W0_clk;
  wire [7:0] mem_121_5_W0_data;
  wire  mem_121_5_W0_en;
  wire  mem_121_5_W0_mask;
  wire [25:0] mem_121_6_R0_addr;
  wire  mem_121_6_R0_clk;
  wire [7:0] mem_121_6_R0_data;
  wire  mem_121_6_R0_en;
  wire [25:0] mem_121_6_W0_addr;
  wire  mem_121_6_W0_clk;
  wire [7:0] mem_121_6_W0_data;
  wire  mem_121_6_W0_en;
  wire  mem_121_6_W0_mask;
  wire [25:0] mem_121_7_R0_addr;
  wire  mem_121_7_R0_clk;
  wire [7:0] mem_121_7_R0_data;
  wire  mem_121_7_R0_en;
  wire [25:0] mem_121_7_W0_addr;
  wire  mem_121_7_W0_clk;
  wire [7:0] mem_121_7_W0_data;
  wire  mem_121_7_W0_en;
  wire  mem_121_7_W0_mask;
  wire [25:0] mem_122_0_R0_addr;
  wire  mem_122_0_R0_clk;
  wire [7:0] mem_122_0_R0_data;
  wire  mem_122_0_R0_en;
  wire [25:0] mem_122_0_W0_addr;
  wire  mem_122_0_W0_clk;
  wire [7:0] mem_122_0_W0_data;
  wire  mem_122_0_W0_en;
  wire  mem_122_0_W0_mask;
  wire [25:0] mem_122_1_R0_addr;
  wire  mem_122_1_R0_clk;
  wire [7:0] mem_122_1_R0_data;
  wire  mem_122_1_R0_en;
  wire [25:0] mem_122_1_W0_addr;
  wire  mem_122_1_W0_clk;
  wire [7:0] mem_122_1_W0_data;
  wire  mem_122_1_W0_en;
  wire  mem_122_1_W0_mask;
  wire [25:0] mem_122_2_R0_addr;
  wire  mem_122_2_R0_clk;
  wire [7:0] mem_122_2_R0_data;
  wire  mem_122_2_R0_en;
  wire [25:0] mem_122_2_W0_addr;
  wire  mem_122_2_W0_clk;
  wire [7:0] mem_122_2_W0_data;
  wire  mem_122_2_W0_en;
  wire  mem_122_2_W0_mask;
  wire [25:0] mem_122_3_R0_addr;
  wire  mem_122_3_R0_clk;
  wire [7:0] mem_122_3_R0_data;
  wire  mem_122_3_R0_en;
  wire [25:0] mem_122_3_W0_addr;
  wire  mem_122_3_W0_clk;
  wire [7:0] mem_122_3_W0_data;
  wire  mem_122_3_W0_en;
  wire  mem_122_3_W0_mask;
  wire [25:0] mem_122_4_R0_addr;
  wire  mem_122_4_R0_clk;
  wire [7:0] mem_122_4_R0_data;
  wire  mem_122_4_R0_en;
  wire [25:0] mem_122_4_W0_addr;
  wire  mem_122_4_W0_clk;
  wire [7:0] mem_122_4_W0_data;
  wire  mem_122_4_W0_en;
  wire  mem_122_4_W0_mask;
  wire [25:0] mem_122_5_R0_addr;
  wire  mem_122_5_R0_clk;
  wire [7:0] mem_122_5_R0_data;
  wire  mem_122_5_R0_en;
  wire [25:0] mem_122_5_W0_addr;
  wire  mem_122_5_W0_clk;
  wire [7:0] mem_122_5_W0_data;
  wire  mem_122_5_W0_en;
  wire  mem_122_5_W0_mask;
  wire [25:0] mem_122_6_R0_addr;
  wire  mem_122_6_R0_clk;
  wire [7:0] mem_122_6_R0_data;
  wire  mem_122_6_R0_en;
  wire [25:0] mem_122_6_W0_addr;
  wire  mem_122_6_W0_clk;
  wire [7:0] mem_122_6_W0_data;
  wire  mem_122_6_W0_en;
  wire  mem_122_6_W0_mask;
  wire [25:0] mem_122_7_R0_addr;
  wire  mem_122_7_R0_clk;
  wire [7:0] mem_122_7_R0_data;
  wire  mem_122_7_R0_en;
  wire [25:0] mem_122_7_W0_addr;
  wire  mem_122_7_W0_clk;
  wire [7:0] mem_122_7_W0_data;
  wire  mem_122_7_W0_en;
  wire  mem_122_7_W0_mask;
  wire [25:0] mem_123_0_R0_addr;
  wire  mem_123_0_R0_clk;
  wire [7:0] mem_123_0_R0_data;
  wire  mem_123_0_R0_en;
  wire [25:0] mem_123_0_W0_addr;
  wire  mem_123_0_W0_clk;
  wire [7:0] mem_123_0_W0_data;
  wire  mem_123_0_W0_en;
  wire  mem_123_0_W0_mask;
  wire [25:0] mem_123_1_R0_addr;
  wire  mem_123_1_R0_clk;
  wire [7:0] mem_123_1_R0_data;
  wire  mem_123_1_R0_en;
  wire [25:0] mem_123_1_W0_addr;
  wire  mem_123_1_W0_clk;
  wire [7:0] mem_123_1_W0_data;
  wire  mem_123_1_W0_en;
  wire  mem_123_1_W0_mask;
  wire [25:0] mem_123_2_R0_addr;
  wire  mem_123_2_R0_clk;
  wire [7:0] mem_123_2_R0_data;
  wire  mem_123_2_R0_en;
  wire [25:0] mem_123_2_W0_addr;
  wire  mem_123_2_W0_clk;
  wire [7:0] mem_123_2_W0_data;
  wire  mem_123_2_W0_en;
  wire  mem_123_2_W0_mask;
  wire [25:0] mem_123_3_R0_addr;
  wire  mem_123_3_R0_clk;
  wire [7:0] mem_123_3_R0_data;
  wire  mem_123_3_R0_en;
  wire [25:0] mem_123_3_W0_addr;
  wire  mem_123_3_W0_clk;
  wire [7:0] mem_123_3_W0_data;
  wire  mem_123_3_W0_en;
  wire  mem_123_3_W0_mask;
  wire [25:0] mem_123_4_R0_addr;
  wire  mem_123_4_R0_clk;
  wire [7:0] mem_123_4_R0_data;
  wire  mem_123_4_R0_en;
  wire [25:0] mem_123_4_W0_addr;
  wire  mem_123_4_W0_clk;
  wire [7:0] mem_123_4_W0_data;
  wire  mem_123_4_W0_en;
  wire  mem_123_4_W0_mask;
  wire [25:0] mem_123_5_R0_addr;
  wire  mem_123_5_R0_clk;
  wire [7:0] mem_123_5_R0_data;
  wire  mem_123_5_R0_en;
  wire [25:0] mem_123_5_W0_addr;
  wire  mem_123_5_W0_clk;
  wire [7:0] mem_123_5_W0_data;
  wire  mem_123_5_W0_en;
  wire  mem_123_5_W0_mask;
  wire [25:0] mem_123_6_R0_addr;
  wire  mem_123_6_R0_clk;
  wire [7:0] mem_123_6_R0_data;
  wire  mem_123_6_R0_en;
  wire [25:0] mem_123_6_W0_addr;
  wire  mem_123_6_W0_clk;
  wire [7:0] mem_123_6_W0_data;
  wire  mem_123_6_W0_en;
  wire  mem_123_6_W0_mask;
  wire [25:0] mem_123_7_R0_addr;
  wire  mem_123_7_R0_clk;
  wire [7:0] mem_123_7_R0_data;
  wire  mem_123_7_R0_en;
  wire [25:0] mem_123_7_W0_addr;
  wire  mem_123_7_W0_clk;
  wire [7:0] mem_123_7_W0_data;
  wire  mem_123_7_W0_en;
  wire  mem_123_7_W0_mask;
  wire [25:0] mem_124_0_R0_addr;
  wire  mem_124_0_R0_clk;
  wire [7:0] mem_124_0_R0_data;
  wire  mem_124_0_R0_en;
  wire [25:0] mem_124_0_W0_addr;
  wire  mem_124_0_W0_clk;
  wire [7:0] mem_124_0_W0_data;
  wire  mem_124_0_W0_en;
  wire  mem_124_0_W0_mask;
  wire [25:0] mem_124_1_R0_addr;
  wire  mem_124_1_R0_clk;
  wire [7:0] mem_124_1_R0_data;
  wire  mem_124_1_R0_en;
  wire [25:0] mem_124_1_W0_addr;
  wire  mem_124_1_W0_clk;
  wire [7:0] mem_124_1_W0_data;
  wire  mem_124_1_W0_en;
  wire  mem_124_1_W0_mask;
  wire [25:0] mem_124_2_R0_addr;
  wire  mem_124_2_R0_clk;
  wire [7:0] mem_124_2_R0_data;
  wire  mem_124_2_R0_en;
  wire [25:0] mem_124_2_W0_addr;
  wire  mem_124_2_W0_clk;
  wire [7:0] mem_124_2_W0_data;
  wire  mem_124_2_W0_en;
  wire  mem_124_2_W0_mask;
  wire [25:0] mem_124_3_R0_addr;
  wire  mem_124_3_R0_clk;
  wire [7:0] mem_124_3_R0_data;
  wire  mem_124_3_R0_en;
  wire [25:0] mem_124_3_W0_addr;
  wire  mem_124_3_W0_clk;
  wire [7:0] mem_124_3_W0_data;
  wire  mem_124_3_W0_en;
  wire  mem_124_3_W0_mask;
  wire [25:0] mem_124_4_R0_addr;
  wire  mem_124_4_R0_clk;
  wire [7:0] mem_124_4_R0_data;
  wire  mem_124_4_R0_en;
  wire [25:0] mem_124_4_W0_addr;
  wire  mem_124_4_W0_clk;
  wire [7:0] mem_124_4_W0_data;
  wire  mem_124_4_W0_en;
  wire  mem_124_4_W0_mask;
  wire [25:0] mem_124_5_R0_addr;
  wire  mem_124_5_R0_clk;
  wire [7:0] mem_124_5_R0_data;
  wire  mem_124_5_R0_en;
  wire [25:0] mem_124_5_W0_addr;
  wire  mem_124_5_W0_clk;
  wire [7:0] mem_124_5_W0_data;
  wire  mem_124_5_W0_en;
  wire  mem_124_5_W0_mask;
  wire [25:0] mem_124_6_R0_addr;
  wire  mem_124_6_R0_clk;
  wire [7:0] mem_124_6_R0_data;
  wire  mem_124_6_R0_en;
  wire [25:0] mem_124_6_W0_addr;
  wire  mem_124_6_W0_clk;
  wire [7:0] mem_124_6_W0_data;
  wire  mem_124_6_W0_en;
  wire  mem_124_6_W0_mask;
  wire [25:0] mem_124_7_R0_addr;
  wire  mem_124_7_R0_clk;
  wire [7:0] mem_124_7_R0_data;
  wire  mem_124_7_R0_en;
  wire [25:0] mem_124_7_W0_addr;
  wire  mem_124_7_W0_clk;
  wire [7:0] mem_124_7_W0_data;
  wire  mem_124_7_W0_en;
  wire  mem_124_7_W0_mask;
  wire [25:0] mem_125_0_R0_addr;
  wire  mem_125_0_R0_clk;
  wire [7:0] mem_125_0_R0_data;
  wire  mem_125_0_R0_en;
  wire [25:0] mem_125_0_W0_addr;
  wire  mem_125_0_W0_clk;
  wire [7:0] mem_125_0_W0_data;
  wire  mem_125_0_W0_en;
  wire  mem_125_0_W0_mask;
  wire [25:0] mem_125_1_R0_addr;
  wire  mem_125_1_R0_clk;
  wire [7:0] mem_125_1_R0_data;
  wire  mem_125_1_R0_en;
  wire [25:0] mem_125_1_W0_addr;
  wire  mem_125_1_W0_clk;
  wire [7:0] mem_125_1_W0_data;
  wire  mem_125_1_W0_en;
  wire  mem_125_1_W0_mask;
  wire [25:0] mem_125_2_R0_addr;
  wire  mem_125_2_R0_clk;
  wire [7:0] mem_125_2_R0_data;
  wire  mem_125_2_R0_en;
  wire [25:0] mem_125_2_W0_addr;
  wire  mem_125_2_W0_clk;
  wire [7:0] mem_125_2_W0_data;
  wire  mem_125_2_W0_en;
  wire  mem_125_2_W0_mask;
  wire [25:0] mem_125_3_R0_addr;
  wire  mem_125_3_R0_clk;
  wire [7:0] mem_125_3_R0_data;
  wire  mem_125_3_R0_en;
  wire [25:0] mem_125_3_W0_addr;
  wire  mem_125_3_W0_clk;
  wire [7:0] mem_125_3_W0_data;
  wire  mem_125_3_W0_en;
  wire  mem_125_3_W0_mask;
  wire [25:0] mem_125_4_R0_addr;
  wire  mem_125_4_R0_clk;
  wire [7:0] mem_125_4_R0_data;
  wire  mem_125_4_R0_en;
  wire [25:0] mem_125_4_W0_addr;
  wire  mem_125_4_W0_clk;
  wire [7:0] mem_125_4_W0_data;
  wire  mem_125_4_W0_en;
  wire  mem_125_4_W0_mask;
  wire [25:0] mem_125_5_R0_addr;
  wire  mem_125_5_R0_clk;
  wire [7:0] mem_125_5_R0_data;
  wire  mem_125_5_R0_en;
  wire [25:0] mem_125_5_W0_addr;
  wire  mem_125_5_W0_clk;
  wire [7:0] mem_125_5_W0_data;
  wire  mem_125_5_W0_en;
  wire  mem_125_5_W0_mask;
  wire [25:0] mem_125_6_R0_addr;
  wire  mem_125_6_R0_clk;
  wire [7:0] mem_125_6_R0_data;
  wire  mem_125_6_R0_en;
  wire [25:0] mem_125_6_W0_addr;
  wire  mem_125_6_W0_clk;
  wire [7:0] mem_125_6_W0_data;
  wire  mem_125_6_W0_en;
  wire  mem_125_6_W0_mask;
  wire [25:0] mem_125_7_R0_addr;
  wire  mem_125_7_R0_clk;
  wire [7:0] mem_125_7_R0_data;
  wire  mem_125_7_R0_en;
  wire [25:0] mem_125_7_W0_addr;
  wire  mem_125_7_W0_clk;
  wire [7:0] mem_125_7_W0_data;
  wire  mem_125_7_W0_en;
  wire  mem_125_7_W0_mask;
  wire [25:0] mem_126_0_R0_addr;
  wire  mem_126_0_R0_clk;
  wire [7:0] mem_126_0_R0_data;
  wire  mem_126_0_R0_en;
  wire [25:0] mem_126_0_W0_addr;
  wire  mem_126_0_W0_clk;
  wire [7:0] mem_126_0_W0_data;
  wire  mem_126_0_W0_en;
  wire  mem_126_0_W0_mask;
  wire [25:0] mem_126_1_R0_addr;
  wire  mem_126_1_R0_clk;
  wire [7:0] mem_126_1_R0_data;
  wire  mem_126_1_R0_en;
  wire [25:0] mem_126_1_W0_addr;
  wire  mem_126_1_W0_clk;
  wire [7:0] mem_126_1_W0_data;
  wire  mem_126_1_W0_en;
  wire  mem_126_1_W0_mask;
  wire [25:0] mem_126_2_R0_addr;
  wire  mem_126_2_R0_clk;
  wire [7:0] mem_126_2_R0_data;
  wire  mem_126_2_R0_en;
  wire [25:0] mem_126_2_W0_addr;
  wire  mem_126_2_W0_clk;
  wire [7:0] mem_126_2_W0_data;
  wire  mem_126_2_W0_en;
  wire  mem_126_2_W0_mask;
  wire [25:0] mem_126_3_R0_addr;
  wire  mem_126_3_R0_clk;
  wire [7:0] mem_126_3_R0_data;
  wire  mem_126_3_R0_en;
  wire [25:0] mem_126_3_W0_addr;
  wire  mem_126_3_W0_clk;
  wire [7:0] mem_126_3_W0_data;
  wire  mem_126_3_W0_en;
  wire  mem_126_3_W0_mask;
  wire [25:0] mem_126_4_R0_addr;
  wire  mem_126_4_R0_clk;
  wire [7:0] mem_126_4_R0_data;
  wire  mem_126_4_R0_en;
  wire [25:0] mem_126_4_W0_addr;
  wire  mem_126_4_W0_clk;
  wire [7:0] mem_126_4_W0_data;
  wire  mem_126_4_W0_en;
  wire  mem_126_4_W0_mask;
  wire [25:0] mem_126_5_R0_addr;
  wire  mem_126_5_R0_clk;
  wire [7:0] mem_126_5_R0_data;
  wire  mem_126_5_R0_en;
  wire [25:0] mem_126_5_W0_addr;
  wire  mem_126_5_W0_clk;
  wire [7:0] mem_126_5_W0_data;
  wire  mem_126_5_W0_en;
  wire  mem_126_5_W0_mask;
  wire [25:0] mem_126_6_R0_addr;
  wire  mem_126_6_R0_clk;
  wire [7:0] mem_126_6_R0_data;
  wire  mem_126_6_R0_en;
  wire [25:0] mem_126_6_W0_addr;
  wire  mem_126_6_W0_clk;
  wire [7:0] mem_126_6_W0_data;
  wire  mem_126_6_W0_en;
  wire  mem_126_6_W0_mask;
  wire [25:0] mem_126_7_R0_addr;
  wire  mem_126_7_R0_clk;
  wire [7:0] mem_126_7_R0_data;
  wire  mem_126_7_R0_en;
  wire [25:0] mem_126_7_W0_addr;
  wire  mem_126_7_W0_clk;
  wire [7:0] mem_126_7_W0_data;
  wire  mem_126_7_W0_en;
  wire  mem_126_7_W0_mask;
  wire [25:0] mem_127_0_R0_addr;
  wire  mem_127_0_R0_clk;
  wire [7:0] mem_127_0_R0_data;
  wire  mem_127_0_R0_en;
  wire [25:0] mem_127_0_W0_addr;
  wire  mem_127_0_W0_clk;
  wire [7:0] mem_127_0_W0_data;
  wire  mem_127_0_W0_en;
  wire  mem_127_0_W0_mask;
  wire [25:0] mem_127_1_R0_addr;
  wire  mem_127_1_R0_clk;
  wire [7:0] mem_127_1_R0_data;
  wire  mem_127_1_R0_en;
  wire [25:0] mem_127_1_W0_addr;
  wire  mem_127_1_W0_clk;
  wire [7:0] mem_127_1_W0_data;
  wire  mem_127_1_W0_en;
  wire  mem_127_1_W0_mask;
  wire [25:0] mem_127_2_R0_addr;
  wire  mem_127_2_R0_clk;
  wire [7:0] mem_127_2_R0_data;
  wire  mem_127_2_R0_en;
  wire [25:0] mem_127_2_W0_addr;
  wire  mem_127_2_W0_clk;
  wire [7:0] mem_127_2_W0_data;
  wire  mem_127_2_W0_en;
  wire  mem_127_2_W0_mask;
  wire [25:0] mem_127_3_R0_addr;
  wire  mem_127_3_R0_clk;
  wire [7:0] mem_127_3_R0_data;
  wire  mem_127_3_R0_en;
  wire [25:0] mem_127_3_W0_addr;
  wire  mem_127_3_W0_clk;
  wire [7:0] mem_127_3_W0_data;
  wire  mem_127_3_W0_en;
  wire  mem_127_3_W0_mask;
  wire [25:0] mem_127_4_R0_addr;
  wire  mem_127_4_R0_clk;
  wire [7:0] mem_127_4_R0_data;
  wire  mem_127_4_R0_en;
  wire [25:0] mem_127_4_W0_addr;
  wire  mem_127_4_W0_clk;
  wire [7:0] mem_127_4_W0_data;
  wire  mem_127_4_W0_en;
  wire  mem_127_4_W0_mask;
  wire [25:0] mem_127_5_R0_addr;
  wire  mem_127_5_R0_clk;
  wire [7:0] mem_127_5_R0_data;
  wire  mem_127_5_R0_en;
  wire [25:0] mem_127_5_W0_addr;
  wire  mem_127_5_W0_clk;
  wire [7:0] mem_127_5_W0_data;
  wire  mem_127_5_W0_en;
  wire  mem_127_5_W0_mask;
  wire [25:0] mem_127_6_R0_addr;
  wire  mem_127_6_R0_clk;
  wire [7:0] mem_127_6_R0_data;
  wire  mem_127_6_R0_en;
  wire [25:0] mem_127_6_W0_addr;
  wire  mem_127_6_W0_clk;
  wire [7:0] mem_127_6_W0_data;
  wire  mem_127_6_W0_en;
  wire  mem_127_6_W0_mask;
  wire [25:0] mem_127_7_R0_addr;
  wire  mem_127_7_R0_clk;
  wire [7:0] mem_127_7_R0_data;
  wire  mem_127_7_R0_en;
  wire [25:0] mem_127_7_W0_addr;
  wire  mem_127_7_W0_clk;
  wire [7:0] mem_127_7_W0_data;
  wire  mem_127_7_W0_en;
  wire  mem_127_7_W0_mask;
  wire [25:0] mem_128_0_R0_addr;
  wire  mem_128_0_R0_clk;
  wire [7:0] mem_128_0_R0_data;
  wire  mem_128_0_R0_en;
  wire [25:0] mem_128_0_W0_addr;
  wire  mem_128_0_W0_clk;
  wire [7:0] mem_128_0_W0_data;
  wire  mem_128_0_W0_en;
  wire  mem_128_0_W0_mask;
  wire [25:0] mem_128_1_R0_addr;
  wire  mem_128_1_R0_clk;
  wire [7:0] mem_128_1_R0_data;
  wire  mem_128_1_R0_en;
  wire [25:0] mem_128_1_W0_addr;
  wire  mem_128_1_W0_clk;
  wire [7:0] mem_128_1_W0_data;
  wire  mem_128_1_W0_en;
  wire  mem_128_1_W0_mask;
  wire [25:0] mem_128_2_R0_addr;
  wire  mem_128_2_R0_clk;
  wire [7:0] mem_128_2_R0_data;
  wire  mem_128_2_R0_en;
  wire [25:0] mem_128_2_W0_addr;
  wire  mem_128_2_W0_clk;
  wire [7:0] mem_128_2_W0_data;
  wire  mem_128_2_W0_en;
  wire  mem_128_2_W0_mask;
  wire [25:0] mem_128_3_R0_addr;
  wire  mem_128_3_R0_clk;
  wire [7:0] mem_128_3_R0_data;
  wire  mem_128_3_R0_en;
  wire [25:0] mem_128_3_W0_addr;
  wire  mem_128_3_W0_clk;
  wire [7:0] mem_128_3_W0_data;
  wire  mem_128_3_W0_en;
  wire  mem_128_3_W0_mask;
  wire [25:0] mem_128_4_R0_addr;
  wire  mem_128_4_R0_clk;
  wire [7:0] mem_128_4_R0_data;
  wire  mem_128_4_R0_en;
  wire [25:0] mem_128_4_W0_addr;
  wire  mem_128_4_W0_clk;
  wire [7:0] mem_128_4_W0_data;
  wire  mem_128_4_W0_en;
  wire  mem_128_4_W0_mask;
  wire [25:0] mem_128_5_R0_addr;
  wire  mem_128_5_R0_clk;
  wire [7:0] mem_128_5_R0_data;
  wire  mem_128_5_R0_en;
  wire [25:0] mem_128_5_W0_addr;
  wire  mem_128_5_W0_clk;
  wire [7:0] mem_128_5_W0_data;
  wire  mem_128_5_W0_en;
  wire  mem_128_5_W0_mask;
  wire [25:0] mem_128_6_R0_addr;
  wire  mem_128_6_R0_clk;
  wire [7:0] mem_128_6_R0_data;
  wire  mem_128_6_R0_en;
  wire [25:0] mem_128_6_W0_addr;
  wire  mem_128_6_W0_clk;
  wire [7:0] mem_128_6_W0_data;
  wire  mem_128_6_W0_en;
  wire  mem_128_6_W0_mask;
  wire [25:0] mem_128_7_R0_addr;
  wire  mem_128_7_R0_clk;
  wire [7:0] mem_128_7_R0_data;
  wire  mem_128_7_R0_en;
  wire [25:0] mem_128_7_W0_addr;
  wire  mem_128_7_W0_clk;
  wire [7:0] mem_128_7_W0_data;
  wire  mem_128_7_W0_en;
  wire  mem_128_7_W0_mask;
  wire [25:0] mem_129_0_R0_addr;
  wire  mem_129_0_R0_clk;
  wire [7:0] mem_129_0_R0_data;
  wire  mem_129_0_R0_en;
  wire [25:0] mem_129_0_W0_addr;
  wire  mem_129_0_W0_clk;
  wire [7:0] mem_129_0_W0_data;
  wire  mem_129_0_W0_en;
  wire  mem_129_0_W0_mask;
  wire [25:0] mem_129_1_R0_addr;
  wire  mem_129_1_R0_clk;
  wire [7:0] mem_129_1_R0_data;
  wire  mem_129_1_R0_en;
  wire [25:0] mem_129_1_W0_addr;
  wire  mem_129_1_W0_clk;
  wire [7:0] mem_129_1_W0_data;
  wire  mem_129_1_W0_en;
  wire  mem_129_1_W0_mask;
  wire [25:0] mem_129_2_R0_addr;
  wire  mem_129_2_R0_clk;
  wire [7:0] mem_129_2_R0_data;
  wire  mem_129_2_R0_en;
  wire [25:0] mem_129_2_W0_addr;
  wire  mem_129_2_W0_clk;
  wire [7:0] mem_129_2_W0_data;
  wire  mem_129_2_W0_en;
  wire  mem_129_2_W0_mask;
  wire [25:0] mem_129_3_R0_addr;
  wire  mem_129_3_R0_clk;
  wire [7:0] mem_129_3_R0_data;
  wire  mem_129_3_R0_en;
  wire [25:0] mem_129_3_W0_addr;
  wire  mem_129_3_W0_clk;
  wire [7:0] mem_129_3_W0_data;
  wire  mem_129_3_W0_en;
  wire  mem_129_3_W0_mask;
  wire [25:0] mem_129_4_R0_addr;
  wire  mem_129_4_R0_clk;
  wire [7:0] mem_129_4_R0_data;
  wire  mem_129_4_R0_en;
  wire [25:0] mem_129_4_W0_addr;
  wire  mem_129_4_W0_clk;
  wire [7:0] mem_129_4_W0_data;
  wire  mem_129_4_W0_en;
  wire  mem_129_4_W0_mask;
  wire [25:0] mem_129_5_R0_addr;
  wire  mem_129_5_R0_clk;
  wire [7:0] mem_129_5_R0_data;
  wire  mem_129_5_R0_en;
  wire [25:0] mem_129_5_W0_addr;
  wire  mem_129_5_W0_clk;
  wire [7:0] mem_129_5_W0_data;
  wire  mem_129_5_W0_en;
  wire  mem_129_5_W0_mask;
  wire [25:0] mem_129_6_R0_addr;
  wire  mem_129_6_R0_clk;
  wire [7:0] mem_129_6_R0_data;
  wire  mem_129_6_R0_en;
  wire [25:0] mem_129_6_W0_addr;
  wire  mem_129_6_W0_clk;
  wire [7:0] mem_129_6_W0_data;
  wire  mem_129_6_W0_en;
  wire  mem_129_6_W0_mask;
  wire [25:0] mem_129_7_R0_addr;
  wire  mem_129_7_R0_clk;
  wire [7:0] mem_129_7_R0_data;
  wire  mem_129_7_R0_en;
  wire [25:0] mem_129_7_W0_addr;
  wire  mem_129_7_W0_clk;
  wire [7:0] mem_129_7_W0_data;
  wire  mem_129_7_W0_en;
  wire  mem_129_7_W0_mask;
  wire [25:0] mem_130_0_R0_addr;
  wire  mem_130_0_R0_clk;
  wire [7:0] mem_130_0_R0_data;
  wire  mem_130_0_R0_en;
  wire [25:0] mem_130_0_W0_addr;
  wire  mem_130_0_W0_clk;
  wire [7:0] mem_130_0_W0_data;
  wire  mem_130_0_W0_en;
  wire  mem_130_0_W0_mask;
  wire [25:0] mem_130_1_R0_addr;
  wire  mem_130_1_R0_clk;
  wire [7:0] mem_130_1_R0_data;
  wire  mem_130_1_R0_en;
  wire [25:0] mem_130_1_W0_addr;
  wire  mem_130_1_W0_clk;
  wire [7:0] mem_130_1_W0_data;
  wire  mem_130_1_W0_en;
  wire  mem_130_1_W0_mask;
  wire [25:0] mem_130_2_R0_addr;
  wire  mem_130_2_R0_clk;
  wire [7:0] mem_130_2_R0_data;
  wire  mem_130_2_R0_en;
  wire [25:0] mem_130_2_W0_addr;
  wire  mem_130_2_W0_clk;
  wire [7:0] mem_130_2_W0_data;
  wire  mem_130_2_W0_en;
  wire  mem_130_2_W0_mask;
  wire [25:0] mem_130_3_R0_addr;
  wire  mem_130_3_R0_clk;
  wire [7:0] mem_130_3_R0_data;
  wire  mem_130_3_R0_en;
  wire [25:0] mem_130_3_W0_addr;
  wire  mem_130_3_W0_clk;
  wire [7:0] mem_130_3_W0_data;
  wire  mem_130_3_W0_en;
  wire  mem_130_3_W0_mask;
  wire [25:0] mem_130_4_R0_addr;
  wire  mem_130_4_R0_clk;
  wire [7:0] mem_130_4_R0_data;
  wire  mem_130_4_R0_en;
  wire [25:0] mem_130_4_W0_addr;
  wire  mem_130_4_W0_clk;
  wire [7:0] mem_130_4_W0_data;
  wire  mem_130_4_W0_en;
  wire  mem_130_4_W0_mask;
  wire [25:0] mem_130_5_R0_addr;
  wire  mem_130_5_R0_clk;
  wire [7:0] mem_130_5_R0_data;
  wire  mem_130_5_R0_en;
  wire [25:0] mem_130_5_W0_addr;
  wire  mem_130_5_W0_clk;
  wire [7:0] mem_130_5_W0_data;
  wire  mem_130_5_W0_en;
  wire  mem_130_5_W0_mask;
  wire [25:0] mem_130_6_R0_addr;
  wire  mem_130_6_R0_clk;
  wire [7:0] mem_130_6_R0_data;
  wire  mem_130_6_R0_en;
  wire [25:0] mem_130_6_W0_addr;
  wire  mem_130_6_W0_clk;
  wire [7:0] mem_130_6_W0_data;
  wire  mem_130_6_W0_en;
  wire  mem_130_6_W0_mask;
  wire [25:0] mem_130_7_R0_addr;
  wire  mem_130_7_R0_clk;
  wire [7:0] mem_130_7_R0_data;
  wire  mem_130_7_R0_en;
  wire [25:0] mem_130_7_W0_addr;
  wire  mem_130_7_W0_clk;
  wire [7:0] mem_130_7_W0_data;
  wire  mem_130_7_W0_en;
  wire  mem_130_7_W0_mask;
  wire [25:0] mem_131_0_R0_addr;
  wire  mem_131_0_R0_clk;
  wire [7:0] mem_131_0_R0_data;
  wire  mem_131_0_R0_en;
  wire [25:0] mem_131_0_W0_addr;
  wire  mem_131_0_W0_clk;
  wire [7:0] mem_131_0_W0_data;
  wire  mem_131_0_W0_en;
  wire  mem_131_0_W0_mask;
  wire [25:0] mem_131_1_R0_addr;
  wire  mem_131_1_R0_clk;
  wire [7:0] mem_131_1_R0_data;
  wire  mem_131_1_R0_en;
  wire [25:0] mem_131_1_W0_addr;
  wire  mem_131_1_W0_clk;
  wire [7:0] mem_131_1_W0_data;
  wire  mem_131_1_W0_en;
  wire  mem_131_1_W0_mask;
  wire [25:0] mem_131_2_R0_addr;
  wire  mem_131_2_R0_clk;
  wire [7:0] mem_131_2_R0_data;
  wire  mem_131_2_R0_en;
  wire [25:0] mem_131_2_W0_addr;
  wire  mem_131_2_W0_clk;
  wire [7:0] mem_131_2_W0_data;
  wire  mem_131_2_W0_en;
  wire  mem_131_2_W0_mask;
  wire [25:0] mem_131_3_R0_addr;
  wire  mem_131_3_R0_clk;
  wire [7:0] mem_131_3_R0_data;
  wire  mem_131_3_R0_en;
  wire [25:0] mem_131_3_W0_addr;
  wire  mem_131_3_W0_clk;
  wire [7:0] mem_131_3_W0_data;
  wire  mem_131_3_W0_en;
  wire  mem_131_3_W0_mask;
  wire [25:0] mem_131_4_R0_addr;
  wire  mem_131_4_R0_clk;
  wire [7:0] mem_131_4_R0_data;
  wire  mem_131_4_R0_en;
  wire [25:0] mem_131_4_W0_addr;
  wire  mem_131_4_W0_clk;
  wire [7:0] mem_131_4_W0_data;
  wire  mem_131_4_W0_en;
  wire  mem_131_4_W0_mask;
  wire [25:0] mem_131_5_R0_addr;
  wire  mem_131_5_R0_clk;
  wire [7:0] mem_131_5_R0_data;
  wire  mem_131_5_R0_en;
  wire [25:0] mem_131_5_W0_addr;
  wire  mem_131_5_W0_clk;
  wire [7:0] mem_131_5_W0_data;
  wire  mem_131_5_W0_en;
  wire  mem_131_5_W0_mask;
  wire [25:0] mem_131_6_R0_addr;
  wire  mem_131_6_R0_clk;
  wire [7:0] mem_131_6_R0_data;
  wire  mem_131_6_R0_en;
  wire [25:0] mem_131_6_W0_addr;
  wire  mem_131_6_W0_clk;
  wire [7:0] mem_131_6_W0_data;
  wire  mem_131_6_W0_en;
  wire  mem_131_6_W0_mask;
  wire [25:0] mem_131_7_R0_addr;
  wire  mem_131_7_R0_clk;
  wire [7:0] mem_131_7_R0_data;
  wire  mem_131_7_R0_en;
  wire [25:0] mem_131_7_W0_addr;
  wire  mem_131_7_W0_clk;
  wire [7:0] mem_131_7_W0_data;
  wire  mem_131_7_W0_en;
  wire  mem_131_7_W0_mask;
  wire [25:0] mem_132_0_R0_addr;
  wire  mem_132_0_R0_clk;
  wire [7:0] mem_132_0_R0_data;
  wire  mem_132_0_R0_en;
  wire [25:0] mem_132_0_W0_addr;
  wire  mem_132_0_W0_clk;
  wire [7:0] mem_132_0_W0_data;
  wire  mem_132_0_W0_en;
  wire  mem_132_0_W0_mask;
  wire [25:0] mem_132_1_R0_addr;
  wire  mem_132_1_R0_clk;
  wire [7:0] mem_132_1_R0_data;
  wire  mem_132_1_R0_en;
  wire [25:0] mem_132_1_W0_addr;
  wire  mem_132_1_W0_clk;
  wire [7:0] mem_132_1_W0_data;
  wire  mem_132_1_W0_en;
  wire  mem_132_1_W0_mask;
  wire [25:0] mem_132_2_R0_addr;
  wire  mem_132_2_R0_clk;
  wire [7:0] mem_132_2_R0_data;
  wire  mem_132_2_R0_en;
  wire [25:0] mem_132_2_W0_addr;
  wire  mem_132_2_W0_clk;
  wire [7:0] mem_132_2_W0_data;
  wire  mem_132_2_W0_en;
  wire  mem_132_2_W0_mask;
  wire [25:0] mem_132_3_R0_addr;
  wire  mem_132_3_R0_clk;
  wire [7:0] mem_132_3_R0_data;
  wire  mem_132_3_R0_en;
  wire [25:0] mem_132_3_W0_addr;
  wire  mem_132_3_W0_clk;
  wire [7:0] mem_132_3_W0_data;
  wire  mem_132_3_W0_en;
  wire  mem_132_3_W0_mask;
  wire [25:0] mem_132_4_R0_addr;
  wire  mem_132_4_R0_clk;
  wire [7:0] mem_132_4_R0_data;
  wire  mem_132_4_R0_en;
  wire [25:0] mem_132_4_W0_addr;
  wire  mem_132_4_W0_clk;
  wire [7:0] mem_132_4_W0_data;
  wire  mem_132_4_W0_en;
  wire  mem_132_4_W0_mask;
  wire [25:0] mem_132_5_R0_addr;
  wire  mem_132_5_R0_clk;
  wire [7:0] mem_132_5_R0_data;
  wire  mem_132_5_R0_en;
  wire [25:0] mem_132_5_W0_addr;
  wire  mem_132_5_W0_clk;
  wire [7:0] mem_132_5_W0_data;
  wire  mem_132_5_W0_en;
  wire  mem_132_5_W0_mask;
  wire [25:0] mem_132_6_R0_addr;
  wire  mem_132_6_R0_clk;
  wire [7:0] mem_132_6_R0_data;
  wire  mem_132_6_R0_en;
  wire [25:0] mem_132_6_W0_addr;
  wire  mem_132_6_W0_clk;
  wire [7:0] mem_132_6_W0_data;
  wire  mem_132_6_W0_en;
  wire  mem_132_6_W0_mask;
  wire [25:0] mem_132_7_R0_addr;
  wire  mem_132_7_R0_clk;
  wire [7:0] mem_132_7_R0_data;
  wire  mem_132_7_R0_en;
  wire [25:0] mem_132_7_W0_addr;
  wire  mem_132_7_W0_clk;
  wire [7:0] mem_132_7_W0_data;
  wire  mem_132_7_W0_en;
  wire  mem_132_7_W0_mask;
  wire [25:0] mem_133_0_R0_addr;
  wire  mem_133_0_R0_clk;
  wire [7:0] mem_133_0_R0_data;
  wire  mem_133_0_R0_en;
  wire [25:0] mem_133_0_W0_addr;
  wire  mem_133_0_W0_clk;
  wire [7:0] mem_133_0_W0_data;
  wire  mem_133_0_W0_en;
  wire  mem_133_0_W0_mask;
  wire [25:0] mem_133_1_R0_addr;
  wire  mem_133_1_R0_clk;
  wire [7:0] mem_133_1_R0_data;
  wire  mem_133_1_R0_en;
  wire [25:0] mem_133_1_W0_addr;
  wire  mem_133_1_W0_clk;
  wire [7:0] mem_133_1_W0_data;
  wire  mem_133_1_W0_en;
  wire  mem_133_1_W0_mask;
  wire [25:0] mem_133_2_R0_addr;
  wire  mem_133_2_R0_clk;
  wire [7:0] mem_133_2_R0_data;
  wire  mem_133_2_R0_en;
  wire [25:0] mem_133_2_W0_addr;
  wire  mem_133_2_W0_clk;
  wire [7:0] mem_133_2_W0_data;
  wire  mem_133_2_W0_en;
  wire  mem_133_2_W0_mask;
  wire [25:0] mem_133_3_R0_addr;
  wire  mem_133_3_R0_clk;
  wire [7:0] mem_133_3_R0_data;
  wire  mem_133_3_R0_en;
  wire [25:0] mem_133_3_W0_addr;
  wire  mem_133_3_W0_clk;
  wire [7:0] mem_133_3_W0_data;
  wire  mem_133_3_W0_en;
  wire  mem_133_3_W0_mask;
  wire [25:0] mem_133_4_R0_addr;
  wire  mem_133_4_R0_clk;
  wire [7:0] mem_133_4_R0_data;
  wire  mem_133_4_R0_en;
  wire [25:0] mem_133_4_W0_addr;
  wire  mem_133_4_W0_clk;
  wire [7:0] mem_133_4_W0_data;
  wire  mem_133_4_W0_en;
  wire  mem_133_4_W0_mask;
  wire [25:0] mem_133_5_R0_addr;
  wire  mem_133_5_R0_clk;
  wire [7:0] mem_133_5_R0_data;
  wire  mem_133_5_R0_en;
  wire [25:0] mem_133_5_W0_addr;
  wire  mem_133_5_W0_clk;
  wire [7:0] mem_133_5_W0_data;
  wire  mem_133_5_W0_en;
  wire  mem_133_5_W0_mask;
  wire [25:0] mem_133_6_R0_addr;
  wire  mem_133_6_R0_clk;
  wire [7:0] mem_133_6_R0_data;
  wire  mem_133_6_R0_en;
  wire [25:0] mem_133_6_W0_addr;
  wire  mem_133_6_W0_clk;
  wire [7:0] mem_133_6_W0_data;
  wire  mem_133_6_W0_en;
  wire  mem_133_6_W0_mask;
  wire [25:0] mem_133_7_R0_addr;
  wire  mem_133_7_R0_clk;
  wire [7:0] mem_133_7_R0_data;
  wire  mem_133_7_R0_en;
  wire [25:0] mem_133_7_W0_addr;
  wire  mem_133_7_W0_clk;
  wire [7:0] mem_133_7_W0_data;
  wire  mem_133_7_W0_en;
  wire  mem_133_7_W0_mask;
  wire [25:0] mem_134_0_R0_addr;
  wire  mem_134_0_R0_clk;
  wire [7:0] mem_134_0_R0_data;
  wire  mem_134_0_R0_en;
  wire [25:0] mem_134_0_W0_addr;
  wire  mem_134_0_W0_clk;
  wire [7:0] mem_134_0_W0_data;
  wire  mem_134_0_W0_en;
  wire  mem_134_0_W0_mask;
  wire [25:0] mem_134_1_R0_addr;
  wire  mem_134_1_R0_clk;
  wire [7:0] mem_134_1_R0_data;
  wire  mem_134_1_R0_en;
  wire [25:0] mem_134_1_W0_addr;
  wire  mem_134_1_W0_clk;
  wire [7:0] mem_134_1_W0_data;
  wire  mem_134_1_W0_en;
  wire  mem_134_1_W0_mask;
  wire [25:0] mem_134_2_R0_addr;
  wire  mem_134_2_R0_clk;
  wire [7:0] mem_134_2_R0_data;
  wire  mem_134_2_R0_en;
  wire [25:0] mem_134_2_W0_addr;
  wire  mem_134_2_W0_clk;
  wire [7:0] mem_134_2_W0_data;
  wire  mem_134_2_W0_en;
  wire  mem_134_2_W0_mask;
  wire [25:0] mem_134_3_R0_addr;
  wire  mem_134_3_R0_clk;
  wire [7:0] mem_134_3_R0_data;
  wire  mem_134_3_R0_en;
  wire [25:0] mem_134_3_W0_addr;
  wire  mem_134_3_W0_clk;
  wire [7:0] mem_134_3_W0_data;
  wire  mem_134_3_W0_en;
  wire  mem_134_3_W0_mask;
  wire [25:0] mem_134_4_R0_addr;
  wire  mem_134_4_R0_clk;
  wire [7:0] mem_134_4_R0_data;
  wire  mem_134_4_R0_en;
  wire [25:0] mem_134_4_W0_addr;
  wire  mem_134_4_W0_clk;
  wire [7:0] mem_134_4_W0_data;
  wire  mem_134_4_W0_en;
  wire  mem_134_4_W0_mask;
  wire [25:0] mem_134_5_R0_addr;
  wire  mem_134_5_R0_clk;
  wire [7:0] mem_134_5_R0_data;
  wire  mem_134_5_R0_en;
  wire [25:0] mem_134_5_W0_addr;
  wire  mem_134_5_W0_clk;
  wire [7:0] mem_134_5_W0_data;
  wire  mem_134_5_W0_en;
  wire  mem_134_5_W0_mask;
  wire [25:0] mem_134_6_R0_addr;
  wire  mem_134_6_R0_clk;
  wire [7:0] mem_134_6_R0_data;
  wire  mem_134_6_R0_en;
  wire [25:0] mem_134_6_W0_addr;
  wire  mem_134_6_W0_clk;
  wire [7:0] mem_134_6_W0_data;
  wire  mem_134_6_W0_en;
  wire  mem_134_6_W0_mask;
  wire [25:0] mem_134_7_R0_addr;
  wire  mem_134_7_R0_clk;
  wire [7:0] mem_134_7_R0_data;
  wire  mem_134_7_R0_en;
  wire [25:0] mem_134_7_W0_addr;
  wire  mem_134_7_W0_clk;
  wire [7:0] mem_134_7_W0_data;
  wire  mem_134_7_W0_en;
  wire  mem_134_7_W0_mask;
  wire [25:0] mem_135_0_R0_addr;
  wire  mem_135_0_R0_clk;
  wire [7:0] mem_135_0_R0_data;
  wire  mem_135_0_R0_en;
  wire [25:0] mem_135_0_W0_addr;
  wire  mem_135_0_W0_clk;
  wire [7:0] mem_135_0_W0_data;
  wire  mem_135_0_W0_en;
  wire  mem_135_0_W0_mask;
  wire [25:0] mem_135_1_R0_addr;
  wire  mem_135_1_R0_clk;
  wire [7:0] mem_135_1_R0_data;
  wire  mem_135_1_R0_en;
  wire [25:0] mem_135_1_W0_addr;
  wire  mem_135_1_W0_clk;
  wire [7:0] mem_135_1_W0_data;
  wire  mem_135_1_W0_en;
  wire  mem_135_1_W0_mask;
  wire [25:0] mem_135_2_R0_addr;
  wire  mem_135_2_R0_clk;
  wire [7:0] mem_135_2_R0_data;
  wire  mem_135_2_R0_en;
  wire [25:0] mem_135_2_W0_addr;
  wire  mem_135_2_W0_clk;
  wire [7:0] mem_135_2_W0_data;
  wire  mem_135_2_W0_en;
  wire  mem_135_2_W0_mask;
  wire [25:0] mem_135_3_R0_addr;
  wire  mem_135_3_R0_clk;
  wire [7:0] mem_135_3_R0_data;
  wire  mem_135_3_R0_en;
  wire [25:0] mem_135_3_W0_addr;
  wire  mem_135_3_W0_clk;
  wire [7:0] mem_135_3_W0_data;
  wire  mem_135_3_W0_en;
  wire  mem_135_3_W0_mask;
  wire [25:0] mem_135_4_R0_addr;
  wire  mem_135_4_R0_clk;
  wire [7:0] mem_135_4_R0_data;
  wire  mem_135_4_R0_en;
  wire [25:0] mem_135_4_W0_addr;
  wire  mem_135_4_W0_clk;
  wire [7:0] mem_135_4_W0_data;
  wire  mem_135_4_W0_en;
  wire  mem_135_4_W0_mask;
  wire [25:0] mem_135_5_R0_addr;
  wire  mem_135_5_R0_clk;
  wire [7:0] mem_135_5_R0_data;
  wire  mem_135_5_R0_en;
  wire [25:0] mem_135_5_W0_addr;
  wire  mem_135_5_W0_clk;
  wire [7:0] mem_135_5_W0_data;
  wire  mem_135_5_W0_en;
  wire  mem_135_5_W0_mask;
  wire [25:0] mem_135_6_R0_addr;
  wire  mem_135_6_R0_clk;
  wire [7:0] mem_135_6_R0_data;
  wire  mem_135_6_R0_en;
  wire [25:0] mem_135_6_W0_addr;
  wire  mem_135_6_W0_clk;
  wire [7:0] mem_135_6_W0_data;
  wire  mem_135_6_W0_en;
  wire  mem_135_6_W0_mask;
  wire [25:0] mem_135_7_R0_addr;
  wire  mem_135_7_R0_clk;
  wire [7:0] mem_135_7_R0_data;
  wire  mem_135_7_R0_en;
  wire [25:0] mem_135_7_W0_addr;
  wire  mem_135_7_W0_clk;
  wire [7:0] mem_135_7_W0_data;
  wire  mem_135_7_W0_en;
  wire  mem_135_7_W0_mask;
  wire [25:0] mem_136_0_R0_addr;
  wire  mem_136_0_R0_clk;
  wire [7:0] mem_136_0_R0_data;
  wire  mem_136_0_R0_en;
  wire [25:0] mem_136_0_W0_addr;
  wire  mem_136_0_W0_clk;
  wire [7:0] mem_136_0_W0_data;
  wire  mem_136_0_W0_en;
  wire  mem_136_0_W0_mask;
  wire [25:0] mem_136_1_R0_addr;
  wire  mem_136_1_R0_clk;
  wire [7:0] mem_136_1_R0_data;
  wire  mem_136_1_R0_en;
  wire [25:0] mem_136_1_W0_addr;
  wire  mem_136_1_W0_clk;
  wire [7:0] mem_136_1_W0_data;
  wire  mem_136_1_W0_en;
  wire  mem_136_1_W0_mask;
  wire [25:0] mem_136_2_R0_addr;
  wire  mem_136_2_R0_clk;
  wire [7:0] mem_136_2_R0_data;
  wire  mem_136_2_R0_en;
  wire [25:0] mem_136_2_W0_addr;
  wire  mem_136_2_W0_clk;
  wire [7:0] mem_136_2_W0_data;
  wire  mem_136_2_W0_en;
  wire  mem_136_2_W0_mask;
  wire [25:0] mem_136_3_R0_addr;
  wire  mem_136_3_R0_clk;
  wire [7:0] mem_136_3_R0_data;
  wire  mem_136_3_R0_en;
  wire [25:0] mem_136_3_W0_addr;
  wire  mem_136_3_W0_clk;
  wire [7:0] mem_136_3_W0_data;
  wire  mem_136_3_W0_en;
  wire  mem_136_3_W0_mask;
  wire [25:0] mem_136_4_R0_addr;
  wire  mem_136_4_R0_clk;
  wire [7:0] mem_136_4_R0_data;
  wire  mem_136_4_R0_en;
  wire [25:0] mem_136_4_W0_addr;
  wire  mem_136_4_W0_clk;
  wire [7:0] mem_136_4_W0_data;
  wire  mem_136_4_W0_en;
  wire  mem_136_4_W0_mask;
  wire [25:0] mem_136_5_R0_addr;
  wire  mem_136_5_R0_clk;
  wire [7:0] mem_136_5_R0_data;
  wire  mem_136_5_R0_en;
  wire [25:0] mem_136_5_W0_addr;
  wire  mem_136_5_W0_clk;
  wire [7:0] mem_136_5_W0_data;
  wire  mem_136_5_W0_en;
  wire  mem_136_5_W0_mask;
  wire [25:0] mem_136_6_R0_addr;
  wire  mem_136_6_R0_clk;
  wire [7:0] mem_136_6_R0_data;
  wire  mem_136_6_R0_en;
  wire [25:0] mem_136_6_W0_addr;
  wire  mem_136_6_W0_clk;
  wire [7:0] mem_136_6_W0_data;
  wire  mem_136_6_W0_en;
  wire  mem_136_6_W0_mask;
  wire [25:0] mem_136_7_R0_addr;
  wire  mem_136_7_R0_clk;
  wire [7:0] mem_136_7_R0_data;
  wire  mem_136_7_R0_en;
  wire [25:0] mem_136_7_W0_addr;
  wire  mem_136_7_W0_clk;
  wire [7:0] mem_136_7_W0_data;
  wire  mem_136_7_W0_en;
  wire  mem_136_7_W0_mask;
  wire [25:0] mem_137_0_R0_addr;
  wire  mem_137_0_R0_clk;
  wire [7:0] mem_137_0_R0_data;
  wire  mem_137_0_R0_en;
  wire [25:0] mem_137_0_W0_addr;
  wire  mem_137_0_W0_clk;
  wire [7:0] mem_137_0_W0_data;
  wire  mem_137_0_W0_en;
  wire  mem_137_0_W0_mask;
  wire [25:0] mem_137_1_R0_addr;
  wire  mem_137_1_R0_clk;
  wire [7:0] mem_137_1_R0_data;
  wire  mem_137_1_R0_en;
  wire [25:0] mem_137_1_W0_addr;
  wire  mem_137_1_W0_clk;
  wire [7:0] mem_137_1_W0_data;
  wire  mem_137_1_W0_en;
  wire  mem_137_1_W0_mask;
  wire [25:0] mem_137_2_R0_addr;
  wire  mem_137_2_R0_clk;
  wire [7:0] mem_137_2_R0_data;
  wire  mem_137_2_R0_en;
  wire [25:0] mem_137_2_W0_addr;
  wire  mem_137_2_W0_clk;
  wire [7:0] mem_137_2_W0_data;
  wire  mem_137_2_W0_en;
  wire  mem_137_2_W0_mask;
  wire [25:0] mem_137_3_R0_addr;
  wire  mem_137_3_R0_clk;
  wire [7:0] mem_137_3_R0_data;
  wire  mem_137_3_R0_en;
  wire [25:0] mem_137_3_W0_addr;
  wire  mem_137_3_W0_clk;
  wire [7:0] mem_137_3_W0_data;
  wire  mem_137_3_W0_en;
  wire  mem_137_3_W0_mask;
  wire [25:0] mem_137_4_R0_addr;
  wire  mem_137_4_R0_clk;
  wire [7:0] mem_137_4_R0_data;
  wire  mem_137_4_R0_en;
  wire [25:0] mem_137_4_W0_addr;
  wire  mem_137_4_W0_clk;
  wire [7:0] mem_137_4_W0_data;
  wire  mem_137_4_W0_en;
  wire  mem_137_4_W0_mask;
  wire [25:0] mem_137_5_R0_addr;
  wire  mem_137_5_R0_clk;
  wire [7:0] mem_137_5_R0_data;
  wire  mem_137_5_R0_en;
  wire [25:0] mem_137_5_W0_addr;
  wire  mem_137_5_W0_clk;
  wire [7:0] mem_137_5_W0_data;
  wire  mem_137_5_W0_en;
  wire  mem_137_5_W0_mask;
  wire [25:0] mem_137_6_R0_addr;
  wire  mem_137_6_R0_clk;
  wire [7:0] mem_137_6_R0_data;
  wire  mem_137_6_R0_en;
  wire [25:0] mem_137_6_W0_addr;
  wire  mem_137_6_W0_clk;
  wire [7:0] mem_137_6_W0_data;
  wire  mem_137_6_W0_en;
  wire  mem_137_6_W0_mask;
  wire [25:0] mem_137_7_R0_addr;
  wire  mem_137_7_R0_clk;
  wire [7:0] mem_137_7_R0_data;
  wire  mem_137_7_R0_en;
  wire [25:0] mem_137_7_W0_addr;
  wire  mem_137_7_W0_clk;
  wire [7:0] mem_137_7_W0_data;
  wire  mem_137_7_W0_en;
  wire  mem_137_7_W0_mask;
  wire [25:0] mem_138_0_R0_addr;
  wire  mem_138_0_R0_clk;
  wire [7:0] mem_138_0_R0_data;
  wire  mem_138_0_R0_en;
  wire [25:0] mem_138_0_W0_addr;
  wire  mem_138_0_W0_clk;
  wire [7:0] mem_138_0_W0_data;
  wire  mem_138_0_W0_en;
  wire  mem_138_0_W0_mask;
  wire [25:0] mem_138_1_R0_addr;
  wire  mem_138_1_R0_clk;
  wire [7:0] mem_138_1_R0_data;
  wire  mem_138_1_R0_en;
  wire [25:0] mem_138_1_W0_addr;
  wire  mem_138_1_W0_clk;
  wire [7:0] mem_138_1_W0_data;
  wire  mem_138_1_W0_en;
  wire  mem_138_1_W0_mask;
  wire [25:0] mem_138_2_R0_addr;
  wire  mem_138_2_R0_clk;
  wire [7:0] mem_138_2_R0_data;
  wire  mem_138_2_R0_en;
  wire [25:0] mem_138_2_W0_addr;
  wire  mem_138_2_W0_clk;
  wire [7:0] mem_138_2_W0_data;
  wire  mem_138_2_W0_en;
  wire  mem_138_2_W0_mask;
  wire [25:0] mem_138_3_R0_addr;
  wire  mem_138_3_R0_clk;
  wire [7:0] mem_138_3_R0_data;
  wire  mem_138_3_R0_en;
  wire [25:0] mem_138_3_W0_addr;
  wire  mem_138_3_W0_clk;
  wire [7:0] mem_138_3_W0_data;
  wire  mem_138_3_W0_en;
  wire  mem_138_3_W0_mask;
  wire [25:0] mem_138_4_R0_addr;
  wire  mem_138_4_R0_clk;
  wire [7:0] mem_138_4_R0_data;
  wire  mem_138_4_R0_en;
  wire [25:0] mem_138_4_W0_addr;
  wire  mem_138_4_W0_clk;
  wire [7:0] mem_138_4_W0_data;
  wire  mem_138_4_W0_en;
  wire  mem_138_4_W0_mask;
  wire [25:0] mem_138_5_R0_addr;
  wire  mem_138_5_R0_clk;
  wire [7:0] mem_138_5_R0_data;
  wire  mem_138_5_R0_en;
  wire [25:0] mem_138_5_W0_addr;
  wire  mem_138_5_W0_clk;
  wire [7:0] mem_138_5_W0_data;
  wire  mem_138_5_W0_en;
  wire  mem_138_5_W0_mask;
  wire [25:0] mem_138_6_R0_addr;
  wire  mem_138_6_R0_clk;
  wire [7:0] mem_138_6_R0_data;
  wire  mem_138_6_R0_en;
  wire [25:0] mem_138_6_W0_addr;
  wire  mem_138_6_W0_clk;
  wire [7:0] mem_138_6_W0_data;
  wire  mem_138_6_W0_en;
  wire  mem_138_6_W0_mask;
  wire [25:0] mem_138_7_R0_addr;
  wire  mem_138_7_R0_clk;
  wire [7:0] mem_138_7_R0_data;
  wire  mem_138_7_R0_en;
  wire [25:0] mem_138_7_W0_addr;
  wire  mem_138_7_W0_clk;
  wire [7:0] mem_138_7_W0_data;
  wire  mem_138_7_W0_en;
  wire  mem_138_7_W0_mask;
  wire [25:0] mem_139_0_R0_addr;
  wire  mem_139_0_R0_clk;
  wire [7:0] mem_139_0_R0_data;
  wire  mem_139_0_R0_en;
  wire [25:0] mem_139_0_W0_addr;
  wire  mem_139_0_W0_clk;
  wire [7:0] mem_139_0_W0_data;
  wire  mem_139_0_W0_en;
  wire  mem_139_0_W0_mask;
  wire [25:0] mem_139_1_R0_addr;
  wire  mem_139_1_R0_clk;
  wire [7:0] mem_139_1_R0_data;
  wire  mem_139_1_R0_en;
  wire [25:0] mem_139_1_W0_addr;
  wire  mem_139_1_W0_clk;
  wire [7:0] mem_139_1_W0_data;
  wire  mem_139_1_W0_en;
  wire  mem_139_1_W0_mask;
  wire [25:0] mem_139_2_R0_addr;
  wire  mem_139_2_R0_clk;
  wire [7:0] mem_139_2_R0_data;
  wire  mem_139_2_R0_en;
  wire [25:0] mem_139_2_W0_addr;
  wire  mem_139_2_W0_clk;
  wire [7:0] mem_139_2_W0_data;
  wire  mem_139_2_W0_en;
  wire  mem_139_2_W0_mask;
  wire [25:0] mem_139_3_R0_addr;
  wire  mem_139_3_R0_clk;
  wire [7:0] mem_139_3_R0_data;
  wire  mem_139_3_R0_en;
  wire [25:0] mem_139_3_W0_addr;
  wire  mem_139_3_W0_clk;
  wire [7:0] mem_139_3_W0_data;
  wire  mem_139_3_W0_en;
  wire  mem_139_3_W0_mask;
  wire [25:0] mem_139_4_R0_addr;
  wire  mem_139_4_R0_clk;
  wire [7:0] mem_139_4_R0_data;
  wire  mem_139_4_R0_en;
  wire [25:0] mem_139_4_W0_addr;
  wire  mem_139_4_W0_clk;
  wire [7:0] mem_139_4_W0_data;
  wire  mem_139_4_W0_en;
  wire  mem_139_4_W0_mask;
  wire [25:0] mem_139_5_R0_addr;
  wire  mem_139_5_R0_clk;
  wire [7:0] mem_139_5_R0_data;
  wire  mem_139_5_R0_en;
  wire [25:0] mem_139_5_W0_addr;
  wire  mem_139_5_W0_clk;
  wire [7:0] mem_139_5_W0_data;
  wire  mem_139_5_W0_en;
  wire  mem_139_5_W0_mask;
  wire [25:0] mem_139_6_R0_addr;
  wire  mem_139_6_R0_clk;
  wire [7:0] mem_139_6_R0_data;
  wire  mem_139_6_R0_en;
  wire [25:0] mem_139_6_W0_addr;
  wire  mem_139_6_W0_clk;
  wire [7:0] mem_139_6_W0_data;
  wire  mem_139_6_W0_en;
  wire  mem_139_6_W0_mask;
  wire [25:0] mem_139_7_R0_addr;
  wire  mem_139_7_R0_clk;
  wire [7:0] mem_139_7_R0_data;
  wire  mem_139_7_R0_en;
  wire [25:0] mem_139_7_W0_addr;
  wire  mem_139_7_W0_clk;
  wire [7:0] mem_139_7_W0_data;
  wire  mem_139_7_W0_en;
  wire  mem_139_7_W0_mask;
  wire [25:0] mem_140_0_R0_addr;
  wire  mem_140_0_R0_clk;
  wire [7:0] mem_140_0_R0_data;
  wire  mem_140_0_R0_en;
  wire [25:0] mem_140_0_W0_addr;
  wire  mem_140_0_W0_clk;
  wire [7:0] mem_140_0_W0_data;
  wire  mem_140_0_W0_en;
  wire  mem_140_0_W0_mask;
  wire [25:0] mem_140_1_R0_addr;
  wire  mem_140_1_R0_clk;
  wire [7:0] mem_140_1_R0_data;
  wire  mem_140_1_R0_en;
  wire [25:0] mem_140_1_W0_addr;
  wire  mem_140_1_W0_clk;
  wire [7:0] mem_140_1_W0_data;
  wire  mem_140_1_W0_en;
  wire  mem_140_1_W0_mask;
  wire [25:0] mem_140_2_R0_addr;
  wire  mem_140_2_R0_clk;
  wire [7:0] mem_140_2_R0_data;
  wire  mem_140_2_R0_en;
  wire [25:0] mem_140_2_W0_addr;
  wire  mem_140_2_W0_clk;
  wire [7:0] mem_140_2_W0_data;
  wire  mem_140_2_W0_en;
  wire  mem_140_2_W0_mask;
  wire [25:0] mem_140_3_R0_addr;
  wire  mem_140_3_R0_clk;
  wire [7:0] mem_140_3_R0_data;
  wire  mem_140_3_R0_en;
  wire [25:0] mem_140_3_W0_addr;
  wire  mem_140_3_W0_clk;
  wire [7:0] mem_140_3_W0_data;
  wire  mem_140_3_W0_en;
  wire  mem_140_3_W0_mask;
  wire [25:0] mem_140_4_R0_addr;
  wire  mem_140_4_R0_clk;
  wire [7:0] mem_140_4_R0_data;
  wire  mem_140_4_R0_en;
  wire [25:0] mem_140_4_W0_addr;
  wire  mem_140_4_W0_clk;
  wire [7:0] mem_140_4_W0_data;
  wire  mem_140_4_W0_en;
  wire  mem_140_4_W0_mask;
  wire [25:0] mem_140_5_R0_addr;
  wire  mem_140_5_R0_clk;
  wire [7:0] mem_140_5_R0_data;
  wire  mem_140_5_R0_en;
  wire [25:0] mem_140_5_W0_addr;
  wire  mem_140_5_W0_clk;
  wire [7:0] mem_140_5_W0_data;
  wire  mem_140_5_W0_en;
  wire  mem_140_5_W0_mask;
  wire [25:0] mem_140_6_R0_addr;
  wire  mem_140_6_R0_clk;
  wire [7:0] mem_140_6_R0_data;
  wire  mem_140_6_R0_en;
  wire [25:0] mem_140_6_W0_addr;
  wire  mem_140_6_W0_clk;
  wire [7:0] mem_140_6_W0_data;
  wire  mem_140_6_W0_en;
  wire  mem_140_6_W0_mask;
  wire [25:0] mem_140_7_R0_addr;
  wire  mem_140_7_R0_clk;
  wire [7:0] mem_140_7_R0_data;
  wire  mem_140_7_R0_en;
  wire [25:0] mem_140_7_W0_addr;
  wire  mem_140_7_W0_clk;
  wire [7:0] mem_140_7_W0_data;
  wire  mem_140_7_W0_en;
  wire  mem_140_7_W0_mask;
  wire [25:0] mem_141_0_R0_addr;
  wire  mem_141_0_R0_clk;
  wire [7:0] mem_141_0_R0_data;
  wire  mem_141_0_R0_en;
  wire [25:0] mem_141_0_W0_addr;
  wire  mem_141_0_W0_clk;
  wire [7:0] mem_141_0_W0_data;
  wire  mem_141_0_W0_en;
  wire  mem_141_0_W0_mask;
  wire [25:0] mem_141_1_R0_addr;
  wire  mem_141_1_R0_clk;
  wire [7:0] mem_141_1_R0_data;
  wire  mem_141_1_R0_en;
  wire [25:0] mem_141_1_W0_addr;
  wire  mem_141_1_W0_clk;
  wire [7:0] mem_141_1_W0_data;
  wire  mem_141_1_W0_en;
  wire  mem_141_1_W0_mask;
  wire [25:0] mem_141_2_R0_addr;
  wire  mem_141_2_R0_clk;
  wire [7:0] mem_141_2_R0_data;
  wire  mem_141_2_R0_en;
  wire [25:0] mem_141_2_W0_addr;
  wire  mem_141_2_W0_clk;
  wire [7:0] mem_141_2_W0_data;
  wire  mem_141_2_W0_en;
  wire  mem_141_2_W0_mask;
  wire [25:0] mem_141_3_R0_addr;
  wire  mem_141_3_R0_clk;
  wire [7:0] mem_141_3_R0_data;
  wire  mem_141_3_R0_en;
  wire [25:0] mem_141_3_W0_addr;
  wire  mem_141_3_W0_clk;
  wire [7:0] mem_141_3_W0_data;
  wire  mem_141_3_W0_en;
  wire  mem_141_3_W0_mask;
  wire [25:0] mem_141_4_R0_addr;
  wire  mem_141_4_R0_clk;
  wire [7:0] mem_141_4_R0_data;
  wire  mem_141_4_R0_en;
  wire [25:0] mem_141_4_W0_addr;
  wire  mem_141_4_W0_clk;
  wire [7:0] mem_141_4_W0_data;
  wire  mem_141_4_W0_en;
  wire  mem_141_4_W0_mask;
  wire [25:0] mem_141_5_R0_addr;
  wire  mem_141_5_R0_clk;
  wire [7:0] mem_141_5_R0_data;
  wire  mem_141_5_R0_en;
  wire [25:0] mem_141_5_W0_addr;
  wire  mem_141_5_W0_clk;
  wire [7:0] mem_141_5_W0_data;
  wire  mem_141_5_W0_en;
  wire  mem_141_5_W0_mask;
  wire [25:0] mem_141_6_R0_addr;
  wire  mem_141_6_R0_clk;
  wire [7:0] mem_141_6_R0_data;
  wire  mem_141_6_R0_en;
  wire [25:0] mem_141_6_W0_addr;
  wire  mem_141_6_W0_clk;
  wire [7:0] mem_141_6_W0_data;
  wire  mem_141_6_W0_en;
  wire  mem_141_6_W0_mask;
  wire [25:0] mem_141_7_R0_addr;
  wire  mem_141_7_R0_clk;
  wire [7:0] mem_141_7_R0_data;
  wire  mem_141_7_R0_en;
  wire [25:0] mem_141_7_W0_addr;
  wire  mem_141_7_W0_clk;
  wire [7:0] mem_141_7_W0_data;
  wire  mem_141_7_W0_en;
  wire  mem_141_7_W0_mask;
  wire [25:0] mem_142_0_R0_addr;
  wire  mem_142_0_R0_clk;
  wire [7:0] mem_142_0_R0_data;
  wire  mem_142_0_R0_en;
  wire [25:0] mem_142_0_W0_addr;
  wire  mem_142_0_W0_clk;
  wire [7:0] mem_142_0_W0_data;
  wire  mem_142_0_W0_en;
  wire  mem_142_0_W0_mask;
  wire [25:0] mem_142_1_R0_addr;
  wire  mem_142_1_R0_clk;
  wire [7:0] mem_142_1_R0_data;
  wire  mem_142_1_R0_en;
  wire [25:0] mem_142_1_W0_addr;
  wire  mem_142_1_W0_clk;
  wire [7:0] mem_142_1_W0_data;
  wire  mem_142_1_W0_en;
  wire  mem_142_1_W0_mask;
  wire [25:0] mem_142_2_R0_addr;
  wire  mem_142_2_R0_clk;
  wire [7:0] mem_142_2_R0_data;
  wire  mem_142_2_R0_en;
  wire [25:0] mem_142_2_W0_addr;
  wire  mem_142_2_W0_clk;
  wire [7:0] mem_142_2_W0_data;
  wire  mem_142_2_W0_en;
  wire  mem_142_2_W0_mask;
  wire [25:0] mem_142_3_R0_addr;
  wire  mem_142_3_R0_clk;
  wire [7:0] mem_142_3_R0_data;
  wire  mem_142_3_R0_en;
  wire [25:0] mem_142_3_W0_addr;
  wire  mem_142_3_W0_clk;
  wire [7:0] mem_142_3_W0_data;
  wire  mem_142_3_W0_en;
  wire  mem_142_3_W0_mask;
  wire [25:0] mem_142_4_R0_addr;
  wire  mem_142_4_R0_clk;
  wire [7:0] mem_142_4_R0_data;
  wire  mem_142_4_R0_en;
  wire [25:0] mem_142_4_W0_addr;
  wire  mem_142_4_W0_clk;
  wire [7:0] mem_142_4_W0_data;
  wire  mem_142_4_W0_en;
  wire  mem_142_4_W0_mask;
  wire [25:0] mem_142_5_R0_addr;
  wire  mem_142_5_R0_clk;
  wire [7:0] mem_142_5_R0_data;
  wire  mem_142_5_R0_en;
  wire [25:0] mem_142_5_W0_addr;
  wire  mem_142_5_W0_clk;
  wire [7:0] mem_142_5_W0_data;
  wire  mem_142_5_W0_en;
  wire  mem_142_5_W0_mask;
  wire [25:0] mem_142_6_R0_addr;
  wire  mem_142_6_R0_clk;
  wire [7:0] mem_142_6_R0_data;
  wire  mem_142_6_R0_en;
  wire [25:0] mem_142_6_W0_addr;
  wire  mem_142_6_W0_clk;
  wire [7:0] mem_142_6_W0_data;
  wire  mem_142_6_W0_en;
  wire  mem_142_6_W0_mask;
  wire [25:0] mem_142_7_R0_addr;
  wire  mem_142_7_R0_clk;
  wire [7:0] mem_142_7_R0_data;
  wire  mem_142_7_R0_en;
  wire [25:0] mem_142_7_W0_addr;
  wire  mem_142_7_W0_clk;
  wire [7:0] mem_142_7_W0_data;
  wire  mem_142_7_W0_en;
  wire  mem_142_7_W0_mask;
  wire [25:0] mem_143_0_R0_addr;
  wire  mem_143_0_R0_clk;
  wire [7:0] mem_143_0_R0_data;
  wire  mem_143_0_R0_en;
  wire [25:0] mem_143_0_W0_addr;
  wire  mem_143_0_W0_clk;
  wire [7:0] mem_143_0_W0_data;
  wire  mem_143_0_W0_en;
  wire  mem_143_0_W0_mask;
  wire [25:0] mem_143_1_R0_addr;
  wire  mem_143_1_R0_clk;
  wire [7:0] mem_143_1_R0_data;
  wire  mem_143_1_R0_en;
  wire [25:0] mem_143_1_W0_addr;
  wire  mem_143_1_W0_clk;
  wire [7:0] mem_143_1_W0_data;
  wire  mem_143_1_W0_en;
  wire  mem_143_1_W0_mask;
  wire [25:0] mem_143_2_R0_addr;
  wire  mem_143_2_R0_clk;
  wire [7:0] mem_143_2_R0_data;
  wire  mem_143_2_R0_en;
  wire [25:0] mem_143_2_W0_addr;
  wire  mem_143_2_W0_clk;
  wire [7:0] mem_143_2_W0_data;
  wire  mem_143_2_W0_en;
  wire  mem_143_2_W0_mask;
  wire [25:0] mem_143_3_R0_addr;
  wire  mem_143_3_R0_clk;
  wire [7:0] mem_143_3_R0_data;
  wire  mem_143_3_R0_en;
  wire [25:0] mem_143_3_W0_addr;
  wire  mem_143_3_W0_clk;
  wire [7:0] mem_143_3_W0_data;
  wire  mem_143_3_W0_en;
  wire  mem_143_3_W0_mask;
  wire [25:0] mem_143_4_R0_addr;
  wire  mem_143_4_R0_clk;
  wire [7:0] mem_143_4_R0_data;
  wire  mem_143_4_R0_en;
  wire [25:0] mem_143_4_W0_addr;
  wire  mem_143_4_W0_clk;
  wire [7:0] mem_143_4_W0_data;
  wire  mem_143_4_W0_en;
  wire  mem_143_4_W0_mask;
  wire [25:0] mem_143_5_R0_addr;
  wire  mem_143_5_R0_clk;
  wire [7:0] mem_143_5_R0_data;
  wire  mem_143_5_R0_en;
  wire [25:0] mem_143_5_W0_addr;
  wire  mem_143_5_W0_clk;
  wire [7:0] mem_143_5_W0_data;
  wire  mem_143_5_W0_en;
  wire  mem_143_5_W0_mask;
  wire [25:0] mem_143_6_R0_addr;
  wire  mem_143_6_R0_clk;
  wire [7:0] mem_143_6_R0_data;
  wire  mem_143_6_R0_en;
  wire [25:0] mem_143_6_W0_addr;
  wire  mem_143_6_W0_clk;
  wire [7:0] mem_143_6_W0_data;
  wire  mem_143_6_W0_en;
  wire  mem_143_6_W0_mask;
  wire [25:0] mem_143_7_R0_addr;
  wire  mem_143_7_R0_clk;
  wire [7:0] mem_143_7_R0_data;
  wire  mem_143_7_R0_en;
  wire [25:0] mem_143_7_W0_addr;
  wire  mem_143_7_W0_clk;
  wire [7:0] mem_143_7_W0_data;
  wire  mem_143_7_W0_en;
  wire  mem_143_7_W0_mask;
  wire [25:0] mem_144_0_R0_addr;
  wire  mem_144_0_R0_clk;
  wire [7:0] mem_144_0_R0_data;
  wire  mem_144_0_R0_en;
  wire [25:0] mem_144_0_W0_addr;
  wire  mem_144_0_W0_clk;
  wire [7:0] mem_144_0_W0_data;
  wire  mem_144_0_W0_en;
  wire  mem_144_0_W0_mask;
  wire [25:0] mem_144_1_R0_addr;
  wire  mem_144_1_R0_clk;
  wire [7:0] mem_144_1_R0_data;
  wire  mem_144_1_R0_en;
  wire [25:0] mem_144_1_W0_addr;
  wire  mem_144_1_W0_clk;
  wire [7:0] mem_144_1_W0_data;
  wire  mem_144_1_W0_en;
  wire  mem_144_1_W0_mask;
  wire [25:0] mem_144_2_R0_addr;
  wire  mem_144_2_R0_clk;
  wire [7:0] mem_144_2_R0_data;
  wire  mem_144_2_R0_en;
  wire [25:0] mem_144_2_W0_addr;
  wire  mem_144_2_W0_clk;
  wire [7:0] mem_144_2_W0_data;
  wire  mem_144_2_W0_en;
  wire  mem_144_2_W0_mask;
  wire [25:0] mem_144_3_R0_addr;
  wire  mem_144_3_R0_clk;
  wire [7:0] mem_144_3_R0_data;
  wire  mem_144_3_R0_en;
  wire [25:0] mem_144_3_W0_addr;
  wire  mem_144_3_W0_clk;
  wire [7:0] mem_144_3_W0_data;
  wire  mem_144_3_W0_en;
  wire  mem_144_3_W0_mask;
  wire [25:0] mem_144_4_R0_addr;
  wire  mem_144_4_R0_clk;
  wire [7:0] mem_144_4_R0_data;
  wire  mem_144_4_R0_en;
  wire [25:0] mem_144_4_W0_addr;
  wire  mem_144_4_W0_clk;
  wire [7:0] mem_144_4_W0_data;
  wire  mem_144_4_W0_en;
  wire  mem_144_4_W0_mask;
  wire [25:0] mem_144_5_R0_addr;
  wire  mem_144_5_R0_clk;
  wire [7:0] mem_144_5_R0_data;
  wire  mem_144_5_R0_en;
  wire [25:0] mem_144_5_W0_addr;
  wire  mem_144_5_W0_clk;
  wire [7:0] mem_144_5_W0_data;
  wire  mem_144_5_W0_en;
  wire  mem_144_5_W0_mask;
  wire [25:0] mem_144_6_R0_addr;
  wire  mem_144_6_R0_clk;
  wire [7:0] mem_144_6_R0_data;
  wire  mem_144_6_R0_en;
  wire [25:0] mem_144_6_W0_addr;
  wire  mem_144_6_W0_clk;
  wire [7:0] mem_144_6_W0_data;
  wire  mem_144_6_W0_en;
  wire  mem_144_6_W0_mask;
  wire [25:0] mem_144_7_R0_addr;
  wire  mem_144_7_R0_clk;
  wire [7:0] mem_144_7_R0_data;
  wire  mem_144_7_R0_en;
  wire [25:0] mem_144_7_W0_addr;
  wire  mem_144_7_W0_clk;
  wire [7:0] mem_144_7_W0_data;
  wire  mem_144_7_W0_en;
  wire  mem_144_7_W0_mask;
  wire [25:0] mem_145_0_R0_addr;
  wire  mem_145_0_R0_clk;
  wire [7:0] mem_145_0_R0_data;
  wire  mem_145_0_R0_en;
  wire [25:0] mem_145_0_W0_addr;
  wire  mem_145_0_W0_clk;
  wire [7:0] mem_145_0_W0_data;
  wire  mem_145_0_W0_en;
  wire  mem_145_0_W0_mask;
  wire [25:0] mem_145_1_R0_addr;
  wire  mem_145_1_R0_clk;
  wire [7:0] mem_145_1_R0_data;
  wire  mem_145_1_R0_en;
  wire [25:0] mem_145_1_W0_addr;
  wire  mem_145_1_W0_clk;
  wire [7:0] mem_145_1_W0_data;
  wire  mem_145_1_W0_en;
  wire  mem_145_1_W0_mask;
  wire [25:0] mem_145_2_R0_addr;
  wire  mem_145_2_R0_clk;
  wire [7:0] mem_145_2_R0_data;
  wire  mem_145_2_R0_en;
  wire [25:0] mem_145_2_W0_addr;
  wire  mem_145_2_W0_clk;
  wire [7:0] mem_145_2_W0_data;
  wire  mem_145_2_W0_en;
  wire  mem_145_2_W0_mask;
  wire [25:0] mem_145_3_R0_addr;
  wire  mem_145_3_R0_clk;
  wire [7:0] mem_145_3_R0_data;
  wire  mem_145_3_R0_en;
  wire [25:0] mem_145_3_W0_addr;
  wire  mem_145_3_W0_clk;
  wire [7:0] mem_145_3_W0_data;
  wire  mem_145_3_W0_en;
  wire  mem_145_3_W0_mask;
  wire [25:0] mem_145_4_R0_addr;
  wire  mem_145_4_R0_clk;
  wire [7:0] mem_145_4_R0_data;
  wire  mem_145_4_R0_en;
  wire [25:0] mem_145_4_W0_addr;
  wire  mem_145_4_W0_clk;
  wire [7:0] mem_145_4_W0_data;
  wire  mem_145_4_W0_en;
  wire  mem_145_4_W0_mask;
  wire [25:0] mem_145_5_R0_addr;
  wire  mem_145_5_R0_clk;
  wire [7:0] mem_145_5_R0_data;
  wire  mem_145_5_R0_en;
  wire [25:0] mem_145_5_W0_addr;
  wire  mem_145_5_W0_clk;
  wire [7:0] mem_145_5_W0_data;
  wire  mem_145_5_W0_en;
  wire  mem_145_5_W0_mask;
  wire [25:0] mem_145_6_R0_addr;
  wire  mem_145_6_R0_clk;
  wire [7:0] mem_145_6_R0_data;
  wire  mem_145_6_R0_en;
  wire [25:0] mem_145_6_W0_addr;
  wire  mem_145_6_W0_clk;
  wire [7:0] mem_145_6_W0_data;
  wire  mem_145_6_W0_en;
  wire  mem_145_6_W0_mask;
  wire [25:0] mem_145_7_R0_addr;
  wire  mem_145_7_R0_clk;
  wire [7:0] mem_145_7_R0_data;
  wire  mem_145_7_R0_en;
  wire [25:0] mem_145_7_W0_addr;
  wire  mem_145_7_W0_clk;
  wire [7:0] mem_145_7_W0_data;
  wire  mem_145_7_W0_en;
  wire  mem_145_7_W0_mask;
  wire [25:0] mem_146_0_R0_addr;
  wire  mem_146_0_R0_clk;
  wire [7:0] mem_146_0_R0_data;
  wire  mem_146_0_R0_en;
  wire [25:0] mem_146_0_W0_addr;
  wire  mem_146_0_W0_clk;
  wire [7:0] mem_146_0_W0_data;
  wire  mem_146_0_W0_en;
  wire  mem_146_0_W0_mask;
  wire [25:0] mem_146_1_R0_addr;
  wire  mem_146_1_R0_clk;
  wire [7:0] mem_146_1_R0_data;
  wire  mem_146_1_R0_en;
  wire [25:0] mem_146_1_W0_addr;
  wire  mem_146_1_W0_clk;
  wire [7:0] mem_146_1_W0_data;
  wire  mem_146_1_W0_en;
  wire  mem_146_1_W0_mask;
  wire [25:0] mem_146_2_R0_addr;
  wire  mem_146_2_R0_clk;
  wire [7:0] mem_146_2_R0_data;
  wire  mem_146_2_R0_en;
  wire [25:0] mem_146_2_W0_addr;
  wire  mem_146_2_W0_clk;
  wire [7:0] mem_146_2_W0_data;
  wire  mem_146_2_W0_en;
  wire  mem_146_2_W0_mask;
  wire [25:0] mem_146_3_R0_addr;
  wire  mem_146_3_R0_clk;
  wire [7:0] mem_146_3_R0_data;
  wire  mem_146_3_R0_en;
  wire [25:0] mem_146_3_W0_addr;
  wire  mem_146_3_W0_clk;
  wire [7:0] mem_146_3_W0_data;
  wire  mem_146_3_W0_en;
  wire  mem_146_3_W0_mask;
  wire [25:0] mem_146_4_R0_addr;
  wire  mem_146_4_R0_clk;
  wire [7:0] mem_146_4_R0_data;
  wire  mem_146_4_R0_en;
  wire [25:0] mem_146_4_W0_addr;
  wire  mem_146_4_W0_clk;
  wire [7:0] mem_146_4_W0_data;
  wire  mem_146_4_W0_en;
  wire  mem_146_4_W0_mask;
  wire [25:0] mem_146_5_R0_addr;
  wire  mem_146_5_R0_clk;
  wire [7:0] mem_146_5_R0_data;
  wire  mem_146_5_R0_en;
  wire [25:0] mem_146_5_W0_addr;
  wire  mem_146_5_W0_clk;
  wire [7:0] mem_146_5_W0_data;
  wire  mem_146_5_W0_en;
  wire  mem_146_5_W0_mask;
  wire [25:0] mem_146_6_R0_addr;
  wire  mem_146_6_R0_clk;
  wire [7:0] mem_146_6_R0_data;
  wire  mem_146_6_R0_en;
  wire [25:0] mem_146_6_W0_addr;
  wire  mem_146_6_W0_clk;
  wire [7:0] mem_146_6_W0_data;
  wire  mem_146_6_W0_en;
  wire  mem_146_6_W0_mask;
  wire [25:0] mem_146_7_R0_addr;
  wire  mem_146_7_R0_clk;
  wire [7:0] mem_146_7_R0_data;
  wire  mem_146_7_R0_en;
  wire [25:0] mem_146_7_W0_addr;
  wire  mem_146_7_W0_clk;
  wire [7:0] mem_146_7_W0_data;
  wire  mem_146_7_W0_en;
  wire  mem_146_7_W0_mask;
  wire [25:0] mem_147_0_R0_addr;
  wire  mem_147_0_R0_clk;
  wire [7:0] mem_147_0_R0_data;
  wire  mem_147_0_R0_en;
  wire [25:0] mem_147_0_W0_addr;
  wire  mem_147_0_W0_clk;
  wire [7:0] mem_147_0_W0_data;
  wire  mem_147_0_W0_en;
  wire  mem_147_0_W0_mask;
  wire [25:0] mem_147_1_R0_addr;
  wire  mem_147_1_R0_clk;
  wire [7:0] mem_147_1_R0_data;
  wire  mem_147_1_R0_en;
  wire [25:0] mem_147_1_W0_addr;
  wire  mem_147_1_W0_clk;
  wire [7:0] mem_147_1_W0_data;
  wire  mem_147_1_W0_en;
  wire  mem_147_1_W0_mask;
  wire [25:0] mem_147_2_R0_addr;
  wire  mem_147_2_R0_clk;
  wire [7:0] mem_147_2_R0_data;
  wire  mem_147_2_R0_en;
  wire [25:0] mem_147_2_W0_addr;
  wire  mem_147_2_W0_clk;
  wire [7:0] mem_147_2_W0_data;
  wire  mem_147_2_W0_en;
  wire  mem_147_2_W0_mask;
  wire [25:0] mem_147_3_R0_addr;
  wire  mem_147_3_R0_clk;
  wire [7:0] mem_147_3_R0_data;
  wire  mem_147_3_R0_en;
  wire [25:0] mem_147_3_W0_addr;
  wire  mem_147_3_W0_clk;
  wire [7:0] mem_147_3_W0_data;
  wire  mem_147_3_W0_en;
  wire  mem_147_3_W0_mask;
  wire [25:0] mem_147_4_R0_addr;
  wire  mem_147_4_R0_clk;
  wire [7:0] mem_147_4_R0_data;
  wire  mem_147_4_R0_en;
  wire [25:0] mem_147_4_W0_addr;
  wire  mem_147_4_W0_clk;
  wire [7:0] mem_147_4_W0_data;
  wire  mem_147_4_W0_en;
  wire  mem_147_4_W0_mask;
  wire [25:0] mem_147_5_R0_addr;
  wire  mem_147_5_R0_clk;
  wire [7:0] mem_147_5_R0_data;
  wire  mem_147_5_R0_en;
  wire [25:0] mem_147_5_W0_addr;
  wire  mem_147_5_W0_clk;
  wire [7:0] mem_147_5_W0_data;
  wire  mem_147_5_W0_en;
  wire  mem_147_5_W0_mask;
  wire [25:0] mem_147_6_R0_addr;
  wire  mem_147_6_R0_clk;
  wire [7:0] mem_147_6_R0_data;
  wire  mem_147_6_R0_en;
  wire [25:0] mem_147_6_W0_addr;
  wire  mem_147_6_W0_clk;
  wire [7:0] mem_147_6_W0_data;
  wire  mem_147_6_W0_en;
  wire  mem_147_6_W0_mask;
  wire [25:0] mem_147_7_R0_addr;
  wire  mem_147_7_R0_clk;
  wire [7:0] mem_147_7_R0_data;
  wire  mem_147_7_R0_en;
  wire [25:0] mem_147_7_W0_addr;
  wire  mem_147_7_W0_clk;
  wire [7:0] mem_147_7_W0_data;
  wire  mem_147_7_W0_en;
  wire  mem_147_7_W0_mask;
  wire [25:0] mem_148_0_R0_addr;
  wire  mem_148_0_R0_clk;
  wire [7:0] mem_148_0_R0_data;
  wire  mem_148_0_R0_en;
  wire [25:0] mem_148_0_W0_addr;
  wire  mem_148_0_W0_clk;
  wire [7:0] mem_148_0_W0_data;
  wire  mem_148_0_W0_en;
  wire  mem_148_0_W0_mask;
  wire [25:0] mem_148_1_R0_addr;
  wire  mem_148_1_R0_clk;
  wire [7:0] mem_148_1_R0_data;
  wire  mem_148_1_R0_en;
  wire [25:0] mem_148_1_W0_addr;
  wire  mem_148_1_W0_clk;
  wire [7:0] mem_148_1_W0_data;
  wire  mem_148_1_W0_en;
  wire  mem_148_1_W0_mask;
  wire [25:0] mem_148_2_R0_addr;
  wire  mem_148_2_R0_clk;
  wire [7:0] mem_148_2_R0_data;
  wire  mem_148_2_R0_en;
  wire [25:0] mem_148_2_W0_addr;
  wire  mem_148_2_W0_clk;
  wire [7:0] mem_148_2_W0_data;
  wire  mem_148_2_W0_en;
  wire  mem_148_2_W0_mask;
  wire [25:0] mem_148_3_R0_addr;
  wire  mem_148_3_R0_clk;
  wire [7:0] mem_148_3_R0_data;
  wire  mem_148_3_R0_en;
  wire [25:0] mem_148_3_W0_addr;
  wire  mem_148_3_W0_clk;
  wire [7:0] mem_148_3_W0_data;
  wire  mem_148_3_W0_en;
  wire  mem_148_3_W0_mask;
  wire [25:0] mem_148_4_R0_addr;
  wire  mem_148_4_R0_clk;
  wire [7:0] mem_148_4_R0_data;
  wire  mem_148_4_R0_en;
  wire [25:0] mem_148_4_W0_addr;
  wire  mem_148_4_W0_clk;
  wire [7:0] mem_148_4_W0_data;
  wire  mem_148_4_W0_en;
  wire  mem_148_4_W0_mask;
  wire [25:0] mem_148_5_R0_addr;
  wire  mem_148_5_R0_clk;
  wire [7:0] mem_148_5_R0_data;
  wire  mem_148_5_R0_en;
  wire [25:0] mem_148_5_W0_addr;
  wire  mem_148_5_W0_clk;
  wire [7:0] mem_148_5_W0_data;
  wire  mem_148_5_W0_en;
  wire  mem_148_5_W0_mask;
  wire [25:0] mem_148_6_R0_addr;
  wire  mem_148_6_R0_clk;
  wire [7:0] mem_148_6_R0_data;
  wire  mem_148_6_R0_en;
  wire [25:0] mem_148_6_W0_addr;
  wire  mem_148_6_W0_clk;
  wire [7:0] mem_148_6_W0_data;
  wire  mem_148_6_W0_en;
  wire  mem_148_6_W0_mask;
  wire [25:0] mem_148_7_R0_addr;
  wire  mem_148_7_R0_clk;
  wire [7:0] mem_148_7_R0_data;
  wire  mem_148_7_R0_en;
  wire [25:0] mem_148_7_W0_addr;
  wire  mem_148_7_W0_clk;
  wire [7:0] mem_148_7_W0_data;
  wire  mem_148_7_W0_en;
  wire  mem_148_7_W0_mask;
  wire [25:0] mem_149_0_R0_addr;
  wire  mem_149_0_R0_clk;
  wire [7:0] mem_149_0_R0_data;
  wire  mem_149_0_R0_en;
  wire [25:0] mem_149_0_W0_addr;
  wire  mem_149_0_W0_clk;
  wire [7:0] mem_149_0_W0_data;
  wire  mem_149_0_W0_en;
  wire  mem_149_0_W0_mask;
  wire [25:0] mem_149_1_R0_addr;
  wire  mem_149_1_R0_clk;
  wire [7:0] mem_149_1_R0_data;
  wire  mem_149_1_R0_en;
  wire [25:0] mem_149_1_W0_addr;
  wire  mem_149_1_W0_clk;
  wire [7:0] mem_149_1_W0_data;
  wire  mem_149_1_W0_en;
  wire  mem_149_1_W0_mask;
  wire [25:0] mem_149_2_R0_addr;
  wire  mem_149_2_R0_clk;
  wire [7:0] mem_149_2_R0_data;
  wire  mem_149_2_R0_en;
  wire [25:0] mem_149_2_W0_addr;
  wire  mem_149_2_W0_clk;
  wire [7:0] mem_149_2_W0_data;
  wire  mem_149_2_W0_en;
  wire  mem_149_2_W0_mask;
  wire [25:0] mem_149_3_R0_addr;
  wire  mem_149_3_R0_clk;
  wire [7:0] mem_149_3_R0_data;
  wire  mem_149_3_R0_en;
  wire [25:0] mem_149_3_W0_addr;
  wire  mem_149_3_W0_clk;
  wire [7:0] mem_149_3_W0_data;
  wire  mem_149_3_W0_en;
  wire  mem_149_3_W0_mask;
  wire [25:0] mem_149_4_R0_addr;
  wire  mem_149_4_R0_clk;
  wire [7:0] mem_149_4_R0_data;
  wire  mem_149_4_R0_en;
  wire [25:0] mem_149_4_W0_addr;
  wire  mem_149_4_W0_clk;
  wire [7:0] mem_149_4_W0_data;
  wire  mem_149_4_W0_en;
  wire  mem_149_4_W0_mask;
  wire [25:0] mem_149_5_R0_addr;
  wire  mem_149_5_R0_clk;
  wire [7:0] mem_149_5_R0_data;
  wire  mem_149_5_R0_en;
  wire [25:0] mem_149_5_W0_addr;
  wire  mem_149_5_W0_clk;
  wire [7:0] mem_149_5_W0_data;
  wire  mem_149_5_W0_en;
  wire  mem_149_5_W0_mask;
  wire [25:0] mem_149_6_R0_addr;
  wire  mem_149_6_R0_clk;
  wire [7:0] mem_149_6_R0_data;
  wire  mem_149_6_R0_en;
  wire [25:0] mem_149_6_W0_addr;
  wire  mem_149_6_W0_clk;
  wire [7:0] mem_149_6_W0_data;
  wire  mem_149_6_W0_en;
  wire  mem_149_6_W0_mask;
  wire [25:0] mem_149_7_R0_addr;
  wire  mem_149_7_R0_clk;
  wire [7:0] mem_149_7_R0_data;
  wire  mem_149_7_R0_en;
  wire [25:0] mem_149_7_W0_addr;
  wire  mem_149_7_W0_clk;
  wire [7:0] mem_149_7_W0_data;
  wire  mem_149_7_W0_en;
  wire  mem_149_7_W0_mask;
  wire [25:0] mem_150_0_R0_addr;
  wire  mem_150_0_R0_clk;
  wire [7:0] mem_150_0_R0_data;
  wire  mem_150_0_R0_en;
  wire [25:0] mem_150_0_W0_addr;
  wire  mem_150_0_W0_clk;
  wire [7:0] mem_150_0_W0_data;
  wire  mem_150_0_W0_en;
  wire  mem_150_0_W0_mask;
  wire [25:0] mem_150_1_R0_addr;
  wire  mem_150_1_R0_clk;
  wire [7:0] mem_150_1_R0_data;
  wire  mem_150_1_R0_en;
  wire [25:0] mem_150_1_W0_addr;
  wire  mem_150_1_W0_clk;
  wire [7:0] mem_150_1_W0_data;
  wire  mem_150_1_W0_en;
  wire  mem_150_1_W0_mask;
  wire [25:0] mem_150_2_R0_addr;
  wire  mem_150_2_R0_clk;
  wire [7:0] mem_150_2_R0_data;
  wire  mem_150_2_R0_en;
  wire [25:0] mem_150_2_W0_addr;
  wire  mem_150_2_W0_clk;
  wire [7:0] mem_150_2_W0_data;
  wire  mem_150_2_W0_en;
  wire  mem_150_2_W0_mask;
  wire [25:0] mem_150_3_R0_addr;
  wire  mem_150_3_R0_clk;
  wire [7:0] mem_150_3_R0_data;
  wire  mem_150_3_R0_en;
  wire [25:0] mem_150_3_W0_addr;
  wire  mem_150_3_W0_clk;
  wire [7:0] mem_150_3_W0_data;
  wire  mem_150_3_W0_en;
  wire  mem_150_3_W0_mask;
  wire [25:0] mem_150_4_R0_addr;
  wire  mem_150_4_R0_clk;
  wire [7:0] mem_150_4_R0_data;
  wire  mem_150_4_R0_en;
  wire [25:0] mem_150_4_W0_addr;
  wire  mem_150_4_W0_clk;
  wire [7:0] mem_150_4_W0_data;
  wire  mem_150_4_W0_en;
  wire  mem_150_4_W0_mask;
  wire [25:0] mem_150_5_R0_addr;
  wire  mem_150_5_R0_clk;
  wire [7:0] mem_150_5_R0_data;
  wire  mem_150_5_R0_en;
  wire [25:0] mem_150_5_W0_addr;
  wire  mem_150_5_W0_clk;
  wire [7:0] mem_150_5_W0_data;
  wire  mem_150_5_W0_en;
  wire  mem_150_5_W0_mask;
  wire [25:0] mem_150_6_R0_addr;
  wire  mem_150_6_R0_clk;
  wire [7:0] mem_150_6_R0_data;
  wire  mem_150_6_R0_en;
  wire [25:0] mem_150_6_W0_addr;
  wire  mem_150_6_W0_clk;
  wire [7:0] mem_150_6_W0_data;
  wire  mem_150_6_W0_en;
  wire  mem_150_6_W0_mask;
  wire [25:0] mem_150_7_R0_addr;
  wire  mem_150_7_R0_clk;
  wire [7:0] mem_150_7_R0_data;
  wire  mem_150_7_R0_en;
  wire [25:0] mem_150_7_W0_addr;
  wire  mem_150_7_W0_clk;
  wire [7:0] mem_150_7_W0_data;
  wire  mem_150_7_W0_en;
  wire  mem_150_7_W0_mask;
  wire [25:0] mem_151_0_R0_addr;
  wire  mem_151_0_R0_clk;
  wire [7:0] mem_151_0_R0_data;
  wire  mem_151_0_R0_en;
  wire [25:0] mem_151_0_W0_addr;
  wire  mem_151_0_W0_clk;
  wire [7:0] mem_151_0_W0_data;
  wire  mem_151_0_W0_en;
  wire  mem_151_0_W0_mask;
  wire [25:0] mem_151_1_R0_addr;
  wire  mem_151_1_R0_clk;
  wire [7:0] mem_151_1_R0_data;
  wire  mem_151_1_R0_en;
  wire [25:0] mem_151_1_W0_addr;
  wire  mem_151_1_W0_clk;
  wire [7:0] mem_151_1_W0_data;
  wire  mem_151_1_W0_en;
  wire  mem_151_1_W0_mask;
  wire [25:0] mem_151_2_R0_addr;
  wire  mem_151_2_R0_clk;
  wire [7:0] mem_151_2_R0_data;
  wire  mem_151_2_R0_en;
  wire [25:0] mem_151_2_W0_addr;
  wire  mem_151_2_W0_clk;
  wire [7:0] mem_151_2_W0_data;
  wire  mem_151_2_W0_en;
  wire  mem_151_2_W0_mask;
  wire [25:0] mem_151_3_R0_addr;
  wire  mem_151_3_R0_clk;
  wire [7:0] mem_151_3_R0_data;
  wire  mem_151_3_R0_en;
  wire [25:0] mem_151_3_W0_addr;
  wire  mem_151_3_W0_clk;
  wire [7:0] mem_151_3_W0_data;
  wire  mem_151_3_W0_en;
  wire  mem_151_3_W0_mask;
  wire [25:0] mem_151_4_R0_addr;
  wire  mem_151_4_R0_clk;
  wire [7:0] mem_151_4_R0_data;
  wire  mem_151_4_R0_en;
  wire [25:0] mem_151_4_W0_addr;
  wire  mem_151_4_W0_clk;
  wire [7:0] mem_151_4_W0_data;
  wire  mem_151_4_W0_en;
  wire  mem_151_4_W0_mask;
  wire [25:0] mem_151_5_R0_addr;
  wire  mem_151_5_R0_clk;
  wire [7:0] mem_151_5_R0_data;
  wire  mem_151_5_R0_en;
  wire [25:0] mem_151_5_W0_addr;
  wire  mem_151_5_W0_clk;
  wire [7:0] mem_151_5_W0_data;
  wire  mem_151_5_W0_en;
  wire  mem_151_5_W0_mask;
  wire [25:0] mem_151_6_R0_addr;
  wire  mem_151_6_R0_clk;
  wire [7:0] mem_151_6_R0_data;
  wire  mem_151_6_R0_en;
  wire [25:0] mem_151_6_W0_addr;
  wire  mem_151_6_W0_clk;
  wire [7:0] mem_151_6_W0_data;
  wire  mem_151_6_W0_en;
  wire  mem_151_6_W0_mask;
  wire [25:0] mem_151_7_R0_addr;
  wire  mem_151_7_R0_clk;
  wire [7:0] mem_151_7_R0_data;
  wire  mem_151_7_R0_en;
  wire [25:0] mem_151_7_W0_addr;
  wire  mem_151_7_W0_clk;
  wire [7:0] mem_151_7_W0_data;
  wire  mem_151_7_W0_en;
  wire  mem_151_7_W0_mask;
  wire [25:0] mem_152_0_R0_addr;
  wire  mem_152_0_R0_clk;
  wire [7:0] mem_152_0_R0_data;
  wire  mem_152_0_R0_en;
  wire [25:0] mem_152_0_W0_addr;
  wire  mem_152_0_W0_clk;
  wire [7:0] mem_152_0_W0_data;
  wire  mem_152_0_W0_en;
  wire  mem_152_0_W0_mask;
  wire [25:0] mem_152_1_R0_addr;
  wire  mem_152_1_R0_clk;
  wire [7:0] mem_152_1_R0_data;
  wire  mem_152_1_R0_en;
  wire [25:0] mem_152_1_W0_addr;
  wire  mem_152_1_W0_clk;
  wire [7:0] mem_152_1_W0_data;
  wire  mem_152_1_W0_en;
  wire  mem_152_1_W0_mask;
  wire [25:0] mem_152_2_R0_addr;
  wire  mem_152_2_R0_clk;
  wire [7:0] mem_152_2_R0_data;
  wire  mem_152_2_R0_en;
  wire [25:0] mem_152_2_W0_addr;
  wire  mem_152_2_W0_clk;
  wire [7:0] mem_152_2_W0_data;
  wire  mem_152_2_W0_en;
  wire  mem_152_2_W0_mask;
  wire [25:0] mem_152_3_R0_addr;
  wire  mem_152_3_R0_clk;
  wire [7:0] mem_152_3_R0_data;
  wire  mem_152_3_R0_en;
  wire [25:0] mem_152_3_W0_addr;
  wire  mem_152_3_W0_clk;
  wire [7:0] mem_152_3_W0_data;
  wire  mem_152_3_W0_en;
  wire  mem_152_3_W0_mask;
  wire [25:0] mem_152_4_R0_addr;
  wire  mem_152_4_R0_clk;
  wire [7:0] mem_152_4_R0_data;
  wire  mem_152_4_R0_en;
  wire [25:0] mem_152_4_W0_addr;
  wire  mem_152_4_W0_clk;
  wire [7:0] mem_152_4_W0_data;
  wire  mem_152_4_W0_en;
  wire  mem_152_4_W0_mask;
  wire [25:0] mem_152_5_R0_addr;
  wire  mem_152_5_R0_clk;
  wire [7:0] mem_152_5_R0_data;
  wire  mem_152_5_R0_en;
  wire [25:0] mem_152_5_W0_addr;
  wire  mem_152_5_W0_clk;
  wire [7:0] mem_152_5_W0_data;
  wire  mem_152_5_W0_en;
  wire  mem_152_5_W0_mask;
  wire [25:0] mem_152_6_R0_addr;
  wire  mem_152_6_R0_clk;
  wire [7:0] mem_152_6_R0_data;
  wire  mem_152_6_R0_en;
  wire [25:0] mem_152_6_W0_addr;
  wire  mem_152_6_W0_clk;
  wire [7:0] mem_152_6_W0_data;
  wire  mem_152_6_W0_en;
  wire  mem_152_6_W0_mask;
  wire [25:0] mem_152_7_R0_addr;
  wire  mem_152_7_R0_clk;
  wire [7:0] mem_152_7_R0_data;
  wire  mem_152_7_R0_en;
  wire [25:0] mem_152_7_W0_addr;
  wire  mem_152_7_W0_clk;
  wire [7:0] mem_152_7_W0_data;
  wire  mem_152_7_W0_en;
  wire  mem_152_7_W0_mask;
  wire [25:0] mem_153_0_R0_addr;
  wire  mem_153_0_R0_clk;
  wire [7:0] mem_153_0_R0_data;
  wire  mem_153_0_R0_en;
  wire [25:0] mem_153_0_W0_addr;
  wire  mem_153_0_W0_clk;
  wire [7:0] mem_153_0_W0_data;
  wire  mem_153_0_W0_en;
  wire  mem_153_0_W0_mask;
  wire [25:0] mem_153_1_R0_addr;
  wire  mem_153_1_R0_clk;
  wire [7:0] mem_153_1_R0_data;
  wire  mem_153_1_R0_en;
  wire [25:0] mem_153_1_W0_addr;
  wire  mem_153_1_W0_clk;
  wire [7:0] mem_153_1_W0_data;
  wire  mem_153_1_W0_en;
  wire  mem_153_1_W0_mask;
  wire [25:0] mem_153_2_R0_addr;
  wire  mem_153_2_R0_clk;
  wire [7:0] mem_153_2_R0_data;
  wire  mem_153_2_R0_en;
  wire [25:0] mem_153_2_W0_addr;
  wire  mem_153_2_W0_clk;
  wire [7:0] mem_153_2_W0_data;
  wire  mem_153_2_W0_en;
  wire  mem_153_2_W0_mask;
  wire [25:0] mem_153_3_R0_addr;
  wire  mem_153_3_R0_clk;
  wire [7:0] mem_153_3_R0_data;
  wire  mem_153_3_R0_en;
  wire [25:0] mem_153_3_W0_addr;
  wire  mem_153_3_W0_clk;
  wire [7:0] mem_153_3_W0_data;
  wire  mem_153_3_W0_en;
  wire  mem_153_3_W0_mask;
  wire [25:0] mem_153_4_R0_addr;
  wire  mem_153_4_R0_clk;
  wire [7:0] mem_153_4_R0_data;
  wire  mem_153_4_R0_en;
  wire [25:0] mem_153_4_W0_addr;
  wire  mem_153_4_W0_clk;
  wire [7:0] mem_153_4_W0_data;
  wire  mem_153_4_W0_en;
  wire  mem_153_4_W0_mask;
  wire [25:0] mem_153_5_R0_addr;
  wire  mem_153_5_R0_clk;
  wire [7:0] mem_153_5_R0_data;
  wire  mem_153_5_R0_en;
  wire [25:0] mem_153_5_W0_addr;
  wire  mem_153_5_W0_clk;
  wire [7:0] mem_153_5_W0_data;
  wire  mem_153_5_W0_en;
  wire  mem_153_5_W0_mask;
  wire [25:0] mem_153_6_R0_addr;
  wire  mem_153_6_R0_clk;
  wire [7:0] mem_153_6_R0_data;
  wire  mem_153_6_R0_en;
  wire [25:0] mem_153_6_W0_addr;
  wire  mem_153_6_W0_clk;
  wire [7:0] mem_153_6_W0_data;
  wire  mem_153_6_W0_en;
  wire  mem_153_6_W0_mask;
  wire [25:0] mem_153_7_R0_addr;
  wire  mem_153_7_R0_clk;
  wire [7:0] mem_153_7_R0_data;
  wire  mem_153_7_R0_en;
  wire [25:0] mem_153_7_W0_addr;
  wire  mem_153_7_W0_clk;
  wire [7:0] mem_153_7_W0_data;
  wire  mem_153_7_W0_en;
  wire  mem_153_7_W0_mask;
  wire [25:0] mem_154_0_R0_addr;
  wire  mem_154_0_R0_clk;
  wire [7:0] mem_154_0_R0_data;
  wire  mem_154_0_R0_en;
  wire [25:0] mem_154_0_W0_addr;
  wire  mem_154_0_W0_clk;
  wire [7:0] mem_154_0_W0_data;
  wire  mem_154_0_W0_en;
  wire  mem_154_0_W0_mask;
  wire [25:0] mem_154_1_R0_addr;
  wire  mem_154_1_R0_clk;
  wire [7:0] mem_154_1_R0_data;
  wire  mem_154_1_R0_en;
  wire [25:0] mem_154_1_W0_addr;
  wire  mem_154_1_W0_clk;
  wire [7:0] mem_154_1_W0_data;
  wire  mem_154_1_W0_en;
  wire  mem_154_1_W0_mask;
  wire [25:0] mem_154_2_R0_addr;
  wire  mem_154_2_R0_clk;
  wire [7:0] mem_154_2_R0_data;
  wire  mem_154_2_R0_en;
  wire [25:0] mem_154_2_W0_addr;
  wire  mem_154_2_W0_clk;
  wire [7:0] mem_154_2_W0_data;
  wire  mem_154_2_W0_en;
  wire  mem_154_2_W0_mask;
  wire [25:0] mem_154_3_R0_addr;
  wire  mem_154_3_R0_clk;
  wire [7:0] mem_154_3_R0_data;
  wire  mem_154_3_R0_en;
  wire [25:0] mem_154_3_W0_addr;
  wire  mem_154_3_W0_clk;
  wire [7:0] mem_154_3_W0_data;
  wire  mem_154_3_W0_en;
  wire  mem_154_3_W0_mask;
  wire [25:0] mem_154_4_R0_addr;
  wire  mem_154_4_R0_clk;
  wire [7:0] mem_154_4_R0_data;
  wire  mem_154_4_R0_en;
  wire [25:0] mem_154_4_W0_addr;
  wire  mem_154_4_W0_clk;
  wire [7:0] mem_154_4_W0_data;
  wire  mem_154_4_W0_en;
  wire  mem_154_4_W0_mask;
  wire [25:0] mem_154_5_R0_addr;
  wire  mem_154_5_R0_clk;
  wire [7:0] mem_154_5_R0_data;
  wire  mem_154_5_R0_en;
  wire [25:0] mem_154_5_W0_addr;
  wire  mem_154_5_W0_clk;
  wire [7:0] mem_154_5_W0_data;
  wire  mem_154_5_W0_en;
  wire  mem_154_5_W0_mask;
  wire [25:0] mem_154_6_R0_addr;
  wire  mem_154_6_R0_clk;
  wire [7:0] mem_154_6_R0_data;
  wire  mem_154_6_R0_en;
  wire [25:0] mem_154_6_W0_addr;
  wire  mem_154_6_W0_clk;
  wire [7:0] mem_154_6_W0_data;
  wire  mem_154_6_W0_en;
  wire  mem_154_6_W0_mask;
  wire [25:0] mem_154_7_R0_addr;
  wire  mem_154_7_R0_clk;
  wire [7:0] mem_154_7_R0_data;
  wire  mem_154_7_R0_en;
  wire [25:0] mem_154_7_W0_addr;
  wire  mem_154_7_W0_clk;
  wire [7:0] mem_154_7_W0_data;
  wire  mem_154_7_W0_en;
  wire  mem_154_7_W0_mask;
  wire [25:0] mem_155_0_R0_addr;
  wire  mem_155_0_R0_clk;
  wire [7:0] mem_155_0_R0_data;
  wire  mem_155_0_R0_en;
  wire [25:0] mem_155_0_W0_addr;
  wire  mem_155_0_W0_clk;
  wire [7:0] mem_155_0_W0_data;
  wire  mem_155_0_W0_en;
  wire  mem_155_0_W0_mask;
  wire [25:0] mem_155_1_R0_addr;
  wire  mem_155_1_R0_clk;
  wire [7:0] mem_155_1_R0_data;
  wire  mem_155_1_R0_en;
  wire [25:0] mem_155_1_W0_addr;
  wire  mem_155_1_W0_clk;
  wire [7:0] mem_155_1_W0_data;
  wire  mem_155_1_W0_en;
  wire  mem_155_1_W0_mask;
  wire [25:0] mem_155_2_R0_addr;
  wire  mem_155_2_R0_clk;
  wire [7:0] mem_155_2_R0_data;
  wire  mem_155_2_R0_en;
  wire [25:0] mem_155_2_W0_addr;
  wire  mem_155_2_W0_clk;
  wire [7:0] mem_155_2_W0_data;
  wire  mem_155_2_W0_en;
  wire  mem_155_2_W0_mask;
  wire [25:0] mem_155_3_R0_addr;
  wire  mem_155_3_R0_clk;
  wire [7:0] mem_155_3_R0_data;
  wire  mem_155_3_R0_en;
  wire [25:0] mem_155_3_W0_addr;
  wire  mem_155_3_W0_clk;
  wire [7:0] mem_155_3_W0_data;
  wire  mem_155_3_W0_en;
  wire  mem_155_3_W0_mask;
  wire [25:0] mem_155_4_R0_addr;
  wire  mem_155_4_R0_clk;
  wire [7:0] mem_155_4_R0_data;
  wire  mem_155_4_R0_en;
  wire [25:0] mem_155_4_W0_addr;
  wire  mem_155_4_W0_clk;
  wire [7:0] mem_155_4_W0_data;
  wire  mem_155_4_W0_en;
  wire  mem_155_4_W0_mask;
  wire [25:0] mem_155_5_R0_addr;
  wire  mem_155_5_R0_clk;
  wire [7:0] mem_155_5_R0_data;
  wire  mem_155_5_R0_en;
  wire [25:0] mem_155_5_W0_addr;
  wire  mem_155_5_W0_clk;
  wire [7:0] mem_155_5_W0_data;
  wire  mem_155_5_W0_en;
  wire  mem_155_5_W0_mask;
  wire [25:0] mem_155_6_R0_addr;
  wire  mem_155_6_R0_clk;
  wire [7:0] mem_155_6_R0_data;
  wire  mem_155_6_R0_en;
  wire [25:0] mem_155_6_W0_addr;
  wire  mem_155_6_W0_clk;
  wire [7:0] mem_155_6_W0_data;
  wire  mem_155_6_W0_en;
  wire  mem_155_6_W0_mask;
  wire [25:0] mem_155_7_R0_addr;
  wire  mem_155_7_R0_clk;
  wire [7:0] mem_155_7_R0_data;
  wire  mem_155_7_R0_en;
  wire [25:0] mem_155_7_W0_addr;
  wire  mem_155_7_W0_clk;
  wire [7:0] mem_155_7_W0_data;
  wire  mem_155_7_W0_en;
  wire  mem_155_7_W0_mask;
  wire [25:0] mem_156_0_R0_addr;
  wire  mem_156_0_R0_clk;
  wire [7:0] mem_156_0_R0_data;
  wire  mem_156_0_R0_en;
  wire [25:0] mem_156_0_W0_addr;
  wire  mem_156_0_W0_clk;
  wire [7:0] mem_156_0_W0_data;
  wire  mem_156_0_W0_en;
  wire  mem_156_0_W0_mask;
  wire [25:0] mem_156_1_R0_addr;
  wire  mem_156_1_R0_clk;
  wire [7:0] mem_156_1_R0_data;
  wire  mem_156_1_R0_en;
  wire [25:0] mem_156_1_W0_addr;
  wire  mem_156_1_W0_clk;
  wire [7:0] mem_156_1_W0_data;
  wire  mem_156_1_W0_en;
  wire  mem_156_1_W0_mask;
  wire [25:0] mem_156_2_R0_addr;
  wire  mem_156_2_R0_clk;
  wire [7:0] mem_156_2_R0_data;
  wire  mem_156_2_R0_en;
  wire [25:0] mem_156_2_W0_addr;
  wire  mem_156_2_W0_clk;
  wire [7:0] mem_156_2_W0_data;
  wire  mem_156_2_W0_en;
  wire  mem_156_2_W0_mask;
  wire [25:0] mem_156_3_R0_addr;
  wire  mem_156_3_R0_clk;
  wire [7:0] mem_156_3_R0_data;
  wire  mem_156_3_R0_en;
  wire [25:0] mem_156_3_W0_addr;
  wire  mem_156_3_W0_clk;
  wire [7:0] mem_156_3_W0_data;
  wire  mem_156_3_W0_en;
  wire  mem_156_3_W0_mask;
  wire [25:0] mem_156_4_R0_addr;
  wire  mem_156_4_R0_clk;
  wire [7:0] mem_156_4_R0_data;
  wire  mem_156_4_R0_en;
  wire [25:0] mem_156_4_W0_addr;
  wire  mem_156_4_W0_clk;
  wire [7:0] mem_156_4_W0_data;
  wire  mem_156_4_W0_en;
  wire  mem_156_4_W0_mask;
  wire [25:0] mem_156_5_R0_addr;
  wire  mem_156_5_R0_clk;
  wire [7:0] mem_156_5_R0_data;
  wire  mem_156_5_R0_en;
  wire [25:0] mem_156_5_W0_addr;
  wire  mem_156_5_W0_clk;
  wire [7:0] mem_156_5_W0_data;
  wire  mem_156_5_W0_en;
  wire  mem_156_5_W0_mask;
  wire [25:0] mem_156_6_R0_addr;
  wire  mem_156_6_R0_clk;
  wire [7:0] mem_156_6_R0_data;
  wire  mem_156_6_R0_en;
  wire [25:0] mem_156_6_W0_addr;
  wire  mem_156_6_W0_clk;
  wire [7:0] mem_156_6_W0_data;
  wire  mem_156_6_W0_en;
  wire  mem_156_6_W0_mask;
  wire [25:0] mem_156_7_R0_addr;
  wire  mem_156_7_R0_clk;
  wire [7:0] mem_156_7_R0_data;
  wire  mem_156_7_R0_en;
  wire [25:0] mem_156_7_W0_addr;
  wire  mem_156_7_W0_clk;
  wire [7:0] mem_156_7_W0_data;
  wire  mem_156_7_W0_en;
  wire  mem_156_7_W0_mask;
  wire [25:0] mem_157_0_R0_addr;
  wire  mem_157_0_R0_clk;
  wire [7:0] mem_157_0_R0_data;
  wire  mem_157_0_R0_en;
  wire [25:0] mem_157_0_W0_addr;
  wire  mem_157_0_W0_clk;
  wire [7:0] mem_157_0_W0_data;
  wire  mem_157_0_W0_en;
  wire  mem_157_0_W0_mask;
  wire [25:0] mem_157_1_R0_addr;
  wire  mem_157_1_R0_clk;
  wire [7:0] mem_157_1_R0_data;
  wire  mem_157_1_R0_en;
  wire [25:0] mem_157_1_W0_addr;
  wire  mem_157_1_W0_clk;
  wire [7:0] mem_157_1_W0_data;
  wire  mem_157_1_W0_en;
  wire  mem_157_1_W0_mask;
  wire [25:0] mem_157_2_R0_addr;
  wire  mem_157_2_R0_clk;
  wire [7:0] mem_157_2_R0_data;
  wire  mem_157_2_R0_en;
  wire [25:0] mem_157_2_W0_addr;
  wire  mem_157_2_W0_clk;
  wire [7:0] mem_157_2_W0_data;
  wire  mem_157_2_W0_en;
  wire  mem_157_2_W0_mask;
  wire [25:0] mem_157_3_R0_addr;
  wire  mem_157_3_R0_clk;
  wire [7:0] mem_157_3_R0_data;
  wire  mem_157_3_R0_en;
  wire [25:0] mem_157_3_W0_addr;
  wire  mem_157_3_W0_clk;
  wire [7:0] mem_157_3_W0_data;
  wire  mem_157_3_W0_en;
  wire  mem_157_3_W0_mask;
  wire [25:0] mem_157_4_R0_addr;
  wire  mem_157_4_R0_clk;
  wire [7:0] mem_157_4_R0_data;
  wire  mem_157_4_R0_en;
  wire [25:0] mem_157_4_W0_addr;
  wire  mem_157_4_W0_clk;
  wire [7:0] mem_157_4_W0_data;
  wire  mem_157_4_W0_en;
  wire  mem_157_4_W0_mask;
  wire [25:0] mem_157_5_R0_addr;
  wire  mem_157_5_R0_clk;
  wire [7:0] mem_157_5_R0_data;
  wire  mem_157_5_R0_en;
  wire [25:0] mem_157_5_W0_addr;
  wire  mem_157_5_W0_clk;
  wire [7:0] mem_157_5_W0_data;
  wire  mem_157_5_W0_en;
  wire  mem_157_5_W0_mask;
  wire [25:0] mem_157_6_R0_addr;
  wire  mem_157_6_R0_clk;
  wire [7:0] mem_157_6_R0_data;
  wire  mem_157_6_R0_en;
  wire [25:0] mem_157_6_W0_addr;
  wire  mem_157_6_W0_clk;
  wire [7:0] mem_157_6_W0_data;
  wire  mem_157_6_W0_en;
  wire  mem_157_6_W0_mask;
  wire [25:0] mem_157_7_R0_addr;
  wire  mem_157_7_R0_clk;
  wire [7:0] mem_157_7_R0_data;
  wire  mem_157_7_R0_en;
  wire [25:0] mem_157_7_W0_addr;
  wire  mem_157_7_W0_clk;
  wire [7:0] mem_157_7_W0_data;
  wire  mem_157_7_W0_en;
  wire  mem_157_7_W0_mask;
  wire [25:0] mem_158_0_R0_addr;
  wire  mem_158_0_R0_clk;
  wire [7:0] mem_158_0_R0_data;
  wire  mem_158_0_R0_en;
  wire [25:0] mem_158_0_W0_addr;
  wire  mem_158_0_W0_clk;
  wire [7:0] mem_158_0_W0_data;
  wire  mem_158_0_W0_en;
  wire  mem_158_0_W0_mask;
  wire [25:0] mem_158_1_R0_addr;
  wire  mem_158_1_R0_clk;
  wire [7:0] mem_158_1_R0_data;
  wire  mem_158_1_R0_en;
  wire [25:0] mem_158_1_W0_addr;
  wire  mem_158_1_W0_clk;
  wire [7:0] mem_158_1_W0_data;
  wire  mem_158_1_W0_en;
  wire  mem_158_1_W0_mask;
  wire [25:0] mem_158_2_R0_addr;
  wire  mem_158_2_R0_clk;
  wire [7:0] mem_158_2_R0_data;
  wire  mem_158_2_R0_en;
  wire [25:0] mem_158_2_W0_addr;
  wire  mem_158_2_W0_clk;
  wire [7:0] mem_158_2_W0_data;
  wire  mem_158_2_W0_en;
  wire  mem_158_2_W0_mask;
  wire [25:0] mem_158_3_R0_addr;
  wire  mem_158_3_R0_clk;
  wire [7:0] mem_158_3_R0_data;
  wire  mem_158_3_R0_en;
  wire [25:0] mem_158_3_W0_addr;
  wire  mem_158_3_W0_clk;
  wire [7:0] mem_158_3_W0_data;
  wire  mem_158_3_W0_en;
  wire  mem_158_3_W0_mask;
  wire [25:0] mem_158_4_R0_addr;
  wire  mem_158_4_R0_clk;
  wire [7:0] mem_158_4_R0_data;
  wire  mem_158_4_R0_en;
  wire [25:0] mem_158_4_W0_addr;
  wire  mem_158_4_W0_clk;
  wire [7:0] mem_158_4_W0_data;
  wire  mem_158_4_W0_en;
  wire  mem_158_4_W0_mask;
  wire [25:0] mem_158_5_R0_addr;
  wire  mem_158_5_R0_clk;
  wire [7:0] mem_158_5_R0_data;
  wire  mem_158_5_R0_en;
  wire [25:0] mem_158_5_W0_addr;
  wire  mem_158_5_W0_clk;
  wire [7:0] mem_158_5_W0_data;
  wire  mem_158_5_W0_en;
  wire  mem_158_5_W0_mask;
  wire [25:0] mem_158_6_R0_addr;
  wire  mem_158_6_R0_clk;
  wire [7:0] mem_158_6_R0_data;
  wire  mem_158_6_R0_en;
  wire [25:0] mem_158_6_W0_addr;
  wire  mem_158_6_W0_clk;
  wire [7:0] mem_158_6_W0_data;
  wire  mem_158_6_W0_en;
  wire  mem_158_6_W0_mask;
  wire [25:0] mem_158_7_R0_addr;
  wire  mem_158_7_R0_clk;
  wire [7:0] mem_158_7_R0_data;
  wire  mem_158_7_R0_en;
  wire [25:0] mem_158_7_W0_addr;
  wire  mem_158_7_W0_clk;
  wire [7:0] mem_158_7_W0_data;
  wire  mem_158_7_W0_en;
  wire  mem_158_7_W0_mask;
  wire [25:0] mem_159_0_R0_addr;
  wire  mem_159_0_R0_clk;
  wire [7:0] mem_159_0_R0_data;
  wire  mem_159_0_R0_en;
  wire [25:0] mem_159_0_W0_addr;
  wire  mem_159_0_W0_clk;
  wire [7:0] mem_159_0_W0_data;
  wire  mem_159_0_W0_en;
  wire  mem_159_0_W0_mask;
  wire [25:0] mem_159_1_R0_addr;
  wire  mem_159_1_R0_clk;
  wire [7:0] mem_159_1_R0_data;
  wire  mem_159_1_R0_en;
  wire [25:0] mem_159_1_W0_addr;
  wire  mem_159_1_W0_clk;
  wire [7:0] mem_159_1_W0_data;
  wire  mem_159_1_W0_en;
  wire  mem_159_1_W0_mask;
  wire [25:0] mem_159_2_R0_addr;
  wire  mem_159_2_R0_clk;
  wire [7:0] mem_159_2_R0_data;
  wire  mem_159_2_R0_en;
  wire [25:0] mem_159_2_W0_addr;
  wire  mem_159_2_W0_clk;
  wire [7:0] mem_159_2_W0_data;
  wire  mem_159_2_W0_en;
  wire  mem_159_2_W0_mask;
  wire [25:0] mem_159_3_R0_addr;
  wire  mem_159_3_R0_clk;
  wire [7:0] mem_159_3_R0_data;
  wire  mem_159_3_R0_en;
  wire [25:0] mem_159_3_W0_addr;
  wire  mem_159_3_W0_clk;
  wire [7:0] mem_159_3_W0_data;
  wire  mem_159_3_W0_en;
  wire  mem_159_3_W0_mask;
  wire [25:0] mem_159_4_R0_addr;
  wire  mem_159_4_R0_clk;
  wire [7:0] mem_159_4_R0_data;
  wire  mem_159_4_R0_en;
  wire [25:0] mem_159_4_W0_addr;
  wire  mem_159_4_W0_clk;
  wire [7:0] mem_159_4_W0_data;
  wire  mem_159_4_W0_en;
  wire  mem_159_4_W0_mask;
  wire [25:0] mem_159_5_R0_addr;
  wire  mem_159_5_R0_clk;
  wire [7:0] mem_159_5_R0_data;
  wire  mem_159_5_R0_en;
  wire [25:0] mem_159_5_W0_addr;
  wire  mem_159_5_W0_clk;
  wire [7:0] mem_159_5_W0_data;
  wire  mem_159_5_W0_en;
  wire  mem_159_5_W0_mask;
  wire [25:0] mem_159_6_R0_addr;
  wire  mem_159_6_R0_clk;
  wire [7:0] mem_159_6_R0_data;
  wire  mem_159_6_R0_en;
  wire [25:0] mem_159_6_W0_addr;
  wire  mem_159_6_W0_clk;
  wire [7:0] mem_159_6_W0_data;
  wire  mem_159_6_W0_en;
  wire  mem_159_6_W0_mask;
  wire [25:0] mem_159_7_R0_addr;
  wire  mem_159_7_R0_clk;
  wire [7:0] mem_159_7_R0_data;
  wire  mem_159_7_R0_en;
  wire [25:0] mem_159_7_W0_addr;
  wire  mem_159_7_W0_clk;
  wire [7:0] mem_159_7_W0_data;
  wire  mem_159_7_W0_en;
  wire  mem_159_7_W0_mask;
  wire [25:0] mem_160_0_R0_addr;
  wire  mem_160_0_R0_clk;
  wire [7:0] mem_160_0_R0_data;
  wire  mem_160_0_R0_en;
  wire [25:0] mem_160_0_W0_addr;
  wire  mem_160_0_W0_clk;
  wire [7:0] mem_160_0_W0_data;
  wire  mem_160_0_W0_en;
  wire  mem_160_0_W0_mask;
  wire [25:0] mem_160_1_R0_addr;
  wire  mem_160_1_R0_clk;
  wire [7:0] mem_160_1_R0_data;
  wire  mem_160_1_R0_en;
  wire [25:0] mem_160_1_W0_addr;
  wire  mem_160_1_W0_clk;
  wire [7:0] mem_160_1_W0_data;
  wire  mem_160_1_W0_en;
  wire  mem_160_1_W0_mask;
  wire [25:0] mem_160_2_R0_addr;
  wire  mem_160_2_R0_clk;
  wire [7:0] mem_160_2_R0_data;
  wire  mem_160_2_R0_en;
  wire [25:0] mem_160_2_W0_addr;
  wire  mem_160_2_W0_clk;
  wire [7:0] mem_160_2_W0_data;
  wire  mem_160_2_W0_en;
  wire  mem_160_2_W0_mask;
  wire [25:0] mem_160_3_R0_addr;
  wire  mem_160_3_R0_clk;
  wire [7:0] mem_160_3_R0_data;
  wire  mem_160_3_R0_en;
  wire [25:0] mem_160_3_W0_addr;
  wire  mem_160_3_W0_clk;
  wire [7:0] mem_160_3_W0_data;
  wire  mem_160_3_W0_en;
  wire  mem_160_3_W0_mask;
  wire [25:0] mem_160_4_R0_addr;
  wire  mem_160_4_R0_clk;
  wire [7:0] mem_160_4_R0_data;
  wire  mem_160_4_R0_en;
  wire [25:0] mem_160_4_W0_addr;
  wire  mem_160_4_W0_clk;
  wire [7:0] mem_160_4_W0_data;
  wire  mem_160_4_W0_en;
  wire  mem_160_4_W0_mask;
  wire [25:0] mem_160_5_R0_addr;
  wire  mem_160_5_R0_clk;
  wire [7:0] mem_160_5_R0_data;
  wire  mem_160_5_R0_en;
  wire [25:0] mem_160_5_W0_addr;
  wire  mem_160_5_W0_clk;
  wire [7:0] mem_160_5_W0_data;
  wire  mem_160_5_W0_en;
  wire  mem_160_5_W0_mask;
  wire [25:0] mem_160_6_R0_addr;
  wire  mem_160_6_R0_clk;
  wire [7:0] mem_160_6_R0_data;
  wire  mem_160_6_R0_en;
  wire [25:0] mem_160_6_W0_addr;
  wire  mem_160_6_W0_clk;
  wire [7:0] mem_160_6_W0_data;
  wire  mem_160_6_W0_en;
  wire  mem_160_6_W0_mask;
  wire [25:0] mem_160_7_R0_addr;
  wire  mem_160_7_R0_clk;
  wire [7:0] mem_160_7_R0_data;
  wire  mem_160_7_R0_en;
  wire [25:0] mem_160_7_W0_addr;
  wire  mem_160_7_W0_clk;
  wire [7:0] mem_160_7_W0_data;
  wire  mem_160_7_W0_en;
  wire  mem_160_7_W0_mask;
  wire [25:0] mem_161_0_R0_addr;
  wire  mem_161_0_R0_clk;
  wire [7:0] mem_161_0_R0_data;
  wire  mem_161_0_R0_en;
  wire [25:0] mem_161_0_W0_addr;
  wire  mem_161_0_W0_clk;
  wire [7:0] mem_161_0_W0_data;
  wire  mem_161_0_W0_en;
  wire  mem_161_0_W0_mask;
  wire [25:0] mem_161_1_R0_addr;
  wire  mem_161_1_R0_clk;
  wire [7:0] mem_161_1_R0_data;
  wire  mem_161_1_R0_en;
  wire [25:0] mem_161_1_W0_addr;
  wire  mem_161_1_W0_clk;
  wire [7:0] mem_161_1_W0_data;
  wire  mem_161_1_W0_en;
  wire  mem_161_1_W0_mask;
  wire [25:0] mem_161_2_R0_addr;
  wire  mem_161_2_R0_clk;
  wire [7:0] mem_161_2_R0_data;
  wire  mem_161_2_R0_en;
  wire [25:0] mem_161_2_W0_addr;
  wire  mem_161_2_W0_clk;
  wire [7:0] mem_161_2_W0_data;
  wire  mem_161_2_W0_en;
  wire  mem_161_2_W0_mask;
  wire [25:0] mem_161_3_R0_addr;
  wire  mem_161_3_R0_clk;
  wire [7:0] mem_161_3_R0_data;
  wire  mem_161_3_R0_en;
  wire [25:0] mem_161_3_W0_addr;
  wire  mem_161_3_W0_clk;
  wire [7:0] mem_161_3_W0_data;
  wire  mem_161_3_W0_en;
  wire  mem_161_3_W0_mask;
  wire [25:0] mem_161_4_R0_addr;
  wire  mem_161_4_R0_clk;
  wire [7:0] mem_161_4_R0_data;
  wire  mem_161_4_R0_en;
  wire [25:0] mem_161_4_W0_addr;
  wire  mem_161_4_W0_clk;
  wire [7:0] mem_161_4_W0_data;
  wire  mem_161_4_W0_en;
  wire  mem_161_4_W0_mask;
  wire [25:0] mem_161_5_R0_addr;
  wire  mem_161_5_R0_clk;
  wire [7:0] mem_161_5_R0_data;
  wire  mem_161_5_R0_en;
  wire [25:0] mem_161_5_W0_addr;
  wire  mem_161_5_W0_clk;
  wire [7:0] mem_161_5_W0_data;
  wire  mem_161_5_W0_en;
  wire  mem_161_5_W0_mask;
  wire [25:0] mem_161_6_R0_addr;
  wire  mem_161_6_R0_clk;
  wire [7:0] mem_161_6_R0_data;
  wire  mem_161_6_R0_en;
  wire [25:0] mem_161_6_W0_addr;
  wire  mem_161_6_W0_clk;
  wire [7:0] mem_161_6_W0_data;
  wire  mem_161_6_W0_en;
  wire  mem_161_6_W0_mask;
  wire [25:0] mem_161_7_R0_addr;
  wire  mem_161_7_R0_clk;
  wire [7:0] mem_161_7_R0_data;
  wire  mem_161_7_R0_en;
  wire [25:0] mem_161_7_W0_addr;
  wire  mem_161_7_W0_clk;
  wire [7:0] mem_161_7_W0_data;
  wire  mem_161_7_W0_en;
  wire  mem_161_7_W0_mask;
  wire [25:0] mem_162_0_R0_addr;
  wire  mem_162_0_R0_clk;
  wire [7:0] mem_162_0_R0_data;
  wire  mem_162_0_R0_en;
  wire [25:0] mem_162_0_W0_addr;
  wire  mem_162_0_W0_clk;
  wire [7:0] mem_162_0_W0_data;
  wire  mem_162_0_W0_en;
  wire  mem_162_0_W0_mask;
  wire [25:0] mem_162_1_R0_addr;
  wire  mem_162_1_R0_clk;
  wire [7:0] mem_162_1_R0_data;
  wire  mem_162_1_R0_en;
  wire [25:0] mem_162_1_W0_addr;
  wire  mem_162_1_W0_clk;
  wire [7:0] mem_162_1_W0_data;
  wire  mem_162_1_W0_en;
  wire  mem_162_1_W0_mask;
  wire [25:0] mem_162_2_R0_addr;
  wire  mem_162_2_R0_clk;
  wire [7:0] mem_162_2_R0_data;
  wire  mem_162_2_R0_en;
  wire [25:0] mem_162_2_W0_addr;
  wire  mem_162_2_W0_clk;
  wire [7:0] mem_162_2_W0_data;
  wire  mem_162_2_W0_en;
  wire  mem_162_2_W0_mask;
  wire [25:0] mem_162_3_R0_addr;
  wire  mem_162_3_R0_clk;
  wire [7:0] mem_162_3_R0_data;
  wire  mem_162_3_R0_en;
  wire [25:0] mem_162_3_W0_addr;
  wire  mem_162_3_W0_clk;
  wire [7:0] mem_162_3_W0_data;
  wire  mem_162_3_W0_en;
  wire  mem_162_3_W0_mask;
  wire [25:0] mem_162_4_R0_addr;
  wire  mem_162_4_R0_clk;
  wire [7:0] mem_162_4_R0_data;
  wire  mem_162_4_R0_en;
  wire [25:0] mem_162_4_W0_addr;
  wire  mem_162_4_W0_clk;
  wire [7:0] mem_162_4_W0_data;
  wire  mem_162_4_W0_en;
  wire  mem_162_4_W0_mask;
  wire [25:0] mem_162_5_R0_addr;
  wire  mem_162_5_R0_clk;
  wire [7:0] mem_162_5_R0_data;
  wire  mem_162_5_R0_en;
  wire [25:0] mem_162_5_W0_addr;
  wire  mem_162_5_W0_clk;
  wire [7:0] mem_162_5_W0_data;
  wire  mem_162_5_W0_en;
  wire  mem_162_5_W0_mask;
  wire [25:0] mem_162_6_R0_addr;
  wire  mem_162_6_R0_clk;
  wire [7:0] mem_162_6_R0_data;
  wire  mem_162_6_R0_en;
  wire [25:0] mem_162_6_W0_addr;
  wire  mem_162_6_W0_clk;
  wire [7:0] mem_162_6_W0_data;
  wire  mem_162_6_W0_en;
  wire  mem_162_6_W0_mask;
  wire [25:0] mem_162_7_R0_addr;
  wire  mem_162_7_R0_clk;
  wire [7:0] mem_162_7_R0_data;
  wire  mem_162_7_R0_en;
  wire [25:0] mem_162_7_W0_addr;
  wire  mem_162_7_W0_clk;
  wire [7:0] mem_162_7_W0_data;
  wire  mem_162_7_W0_en;
  wire  mem_162_7_W0_mask;
  wire [25:0] mem_163_0_R0_addr;
  wire  mem_163_0_R0_clk;
  wire [7:0] mem_163_0_R0_data;
  wire  mem_163_0_R0_en;
  wire [25:0] mem_163_0_W0_addr;
  wire  mem_163_0_W0_clk;
  wire [7:0] mem_163_0_W0_data;
  wire  mem_163_0_W0_en;
  wire  mem_163_0_W0_mask;
  wire [25:0] mem_163_1_R0_addr;
  wire  mem_163_1_R0_clk;
  wire [7:0] mem_163_1_R0_data;
  wire  mem_163_1_R0_en;
  wire [25:0] mem_163_1_W0_addr;
  wire  mem_163_1_W0_clk;
  wire [7:0] mem_163_1_W0_data;
  wire  mem_163_1_W0_en;
  wire  mem_163_1_W0_mask;
  wire [25:0] mem_163_2_R0_addr;
  wire  mem_163_2_R0_clk;
  wire [7:0] mem_163_2_R0_data;
  wire  mem_163_2_R0_en;
  wire [25:0] mem_163_2_W0_addr;
  wire  mem_163_2_W0_clk;
  wire [7:0] mem_163_2_W0_data;
  wire  mem_163_2_W0_en;
  wire  mem_163_2_W0_mask;
  wire [25:0] mem_163_3_R0_addr;
  wire  mem_163_3_R0_clk;
  wire [7:0] mem_163_3_R0_data;
  wire  mem_163_3_R0_en;
  wire [25:0] mem_163_3_W0_addr;
  wire  mem_163_3_W0_clk;
  wire [7:0] mem_163_3_W0_data;
  wire  mem_163_3_W0_en;
  wire  mem_163_3_W0_mask;
  wire [25:0] mem_163_4_R0_addr;
  wire  mem_163_4_R0_clk;
  wire [7:0] mem_163_4_R0_data;
  wire  mem_163_4_R0_en;
  wire [25:0] mem_163_4_W0_addr;
  wire  mem_163_4_W0_clk;
  wire [7:0] mem_163_4_W0_data;
  wire  mem_163_4_W0_en;
  wire  mem_163_4_W0_mask;
  wire [25:0] mem_163_5_R0_addr;
  wire  mem_163_5_R0_clk;
  wire [7:0] mem_163_5_R0_data;
  wire  mem_163_5_R0_en;
  wire [25:0] mem_163_5_W0_addr;
  wire  mem_163_5_W0_clk;
  wire [7:0] mem_163_5_W0_data;
  wire  mem_163_5_W0_en;
  wire  mem_163_5_W0_mask;
  wire [25:0] mem_163_6_R0_addr;
  wire  mem_163_6_R0_clk;
  wire [7:0] mem_163_6_R0_data;
  wire  mem_163_6_R0_en;
  wire [25:0] mem_163_6_W0_addr;
  wire  mem_163_6_W0_clk;
  wire [7:0] mem_163_6_W0_data;
  wire  mem_163_6_W0_en;
  wire  mem_163_6_W0_mask;
  wire [25:0] mem_163_7_R0_addr;
  wire  mem_163_7_R0_clk;
  wire [7:0] mem_163_7_R0_data;
  wire  mem_163_7_R0_en;
  wire [25:0] mem_163_7_W0_addr;
  wire  mem_163_7_W0_clk;
  wire [7:0] mem_163_7_W0_data;
  wire  mem_163_7_W0_en;
  wire  mem_163_7_W0_mask;
  wire [25:0] mem_164_0_R0_addr;
  wire  mem_164_0_R0_clk;
  wire [7:0] mem_164_0_R0_data;
  wire  mem_164_0_R0_en;
  wire [25:0] mem_164_0_W0_addr;
  wire  mem_164_0_W0_clk;
  wire [7:0] mem_164_0_W0_data;
  wire  mem_164_0_W0_en;
  wire  mem_164_0_W0_mask;
  wire [25:0] mem_164_1_R0_addr;
  wire  mem_164_1_R0_clk;
  wire [7:0] mem_164_1_R0_data;
  wire  mem_164_1_R0_en;
  wire [25:0] mem_164_1_W0_addr;
  wire  mem_164_1_W0_clk;
  wire [7:0] mem_164_1_W0_data;
  wire  mem_164_1_W0_en;
  wire  mem_164_1_W0_mask;
  wire [25:0] mem_164_2_R0_addr;
  wire  mem_164_2_R0_clk;
  wire [7:0] mem_164_2_R0_data;
  wire  mem_164_2_R0_en;
  wire [25:0] mem_164_2_W0_addr;
  wire  mem_164_2_W0_clk;
  wire [7:0] mem_164_2_W0_data;
  wire  mem_164_2_W0_en;
  wire  mem_164_2_W0_mask;
  wire [25:0] mem_164_3_R0_addr;
  wire  mem_164_3_R0_clk;
  wire [7:0] mem_164_3_R0_data;
  wire  mem_164_3_R0_en;
  wire [25:0] mem_164_3_W0_addr;
  wire  mem_164_3_W0_clk;
  wire [7:0] mem_164_3_W0_data;
  wire  mem_164_3_W0_en;
  wire  mem_164_3_W0_mask;
  wire [25:0] mem_164_4_R0_addr;
  wire  mem_164_4_R0_clk;
  wire [7:0] mem_164_4_R0_data;
  wire  mem_164_4_R0_en;
  wire [25:0] mem_164_4_W0_addr;
  wire  mem_164_4_W0_clk;
  wire [7:0] mem_164_4_W0_data;
  wire  mem_164_4_W0_en;
  wire  mem_164_4_W0_mask;
  wire [25:0] mem_164_5_R0_addr;
  wire  mem_164_5_R0_clk;
  wire [7:0] mem_164_5_R0_data;
  wire  mem_164_5_R0_en;
  wire [25:0] mem_164_5_W0_addr;
  wire  mem_164_5_W0_clk;
  wire [7:0] mem_164_5_W0_data;
  wire  mem_164_5_W0_en;
  wire  mem_164_5_W0_mask;
  wire [25:0] mem_164_6_R0_addr;
  wire  mem_164_6_R0_clk;
  wire [7:0] mem_164_6_R0_data;
  wire  mem_164_6_R0_en;
  wire [25:0] mem_164_6_W0_addr;
  wire  mem_164_6_W0_clk;
  wire [7:0] mem_164_6_W0_data;
  wire  mem_164_6_W0_en;
  wire  mem_164_6_W0_mask;
  wire [25:0] mem_164_7_R0_addr;
  wire  mem_164_7_R0_clk;
  wire [7:0] mem_164_7_R0_data;
  wire  mem_164_7_R0_en;
  wire [25:0] mem_164_7_W0_addr;
  wire  mem_164_7_W0_clk;
  wire [7:0] mem_164_7_W0_data;
  wire  mem_164_7_W0_en;
  wire  mem_164_7_W0_mask;
  wire [25:0] mem_165_0_R0_addr;
  wire  mem_165_0_R0_clk;
  wire [7:0] mem_165_0_R0_data;
  wire  mem_165_0_R0_en;
  wire [25:0] mem_165_0_W0_addr;
  wire  mem_165_0_W0_clk;
  wire [7:0] mem_165_0_W0_data;
  wire  mem_165_0_W0_en;
  wire  mem_165_0_W0_mask;
  wire [25:0] mem_165_1_R0_addr;
  wire  mem_165_1_R0_clk;
  wire [7:0] mem_165_1_R0_data;
  wire  mem_165_1_R0_en;
  wire [25:0] mem_165_1_W0_addr;
  wire  mem_165_1_W0_clk;
  wire [7:0] mem_165_1_W0_data;
  wire  mem_165_1_W0_en;
  wire  mem_165_1_W0_mask;
  wire [25:0] mem_165_2_R0_addr;
  wire  mem_165_2_R0_clk;
  wire [7:0] mem_165_2_R0_data;
  wire  mem_165_2_R0_en;
  wire [25:0] mem_165_2_W0_addr;
  wire  mem_165_2_W0_clk;
  wire [7:0] mem_165_2_W0_data;
  wire  mem_165_2_W0_en;
  wire  mem_165_2_W0_mask;
  wire [25:0] mem_165_3_R0_addr;
  wire  mem_165_3_R0_clk;
  wire [7:0] mem_165_3_R0_data;
  wire  mem_165_3_R0_en;
  wire [25:0] mem_165_3_W0_addr;
  wire  mem_165_3_W0_clk;
  wire [7:0] mem_165_3_W0_data;
  wire  mem_165_3_W0_en;
  wire  mem_165_3_W0_mask;
  wire [25:0] mem_165_4_R0_addr;
  wire  mem_165_4_R0_clk;
  wire [7:0] mem_165_4_R0_data;
  wire  mem_165_4_R0_en;
  wire [25:0] mem_165_4_W0_addr;
  wire  mem_165_4_W0_clk;
  wire [7:0] mem_165_4_W0_data;
  wire  mem_165_4_W0_en;
  wire  mem_165_4_W0_mask;
  wire [25:0] mem_165_5_R0_addr;
  wire  mem_165_5_R0_clk;
  wire [7:0] mem_165_5_R0_data;
  wire  mem_165_5_R0_en;
  wire [25:0] mem_165_5_W0_addr;
  wire  mem_165_5_W0_clk;
  wire [7:0] mem_165_5_W0_data;
  wire  mem_165_5_W0_en;
  wire  mem_165_5_W0_mask;
  wire [25:0] mem_165_6_R0_addr;
  wire  mem_165_6_R0_clk;
  wire [7:0] mem_165_6_R0_data;
  wire  mem_165_6_R0_en;
  wire [25:0] mem_165_6_W0_addr;
  wire  mem_165_6_W0_clk;
  wire [7:0] mem_165_6_W0_data;
  wire  mem_165_6_W0_en;
  wire  mem_165_6_W0_mask;
  wire [25:0] mem_165_7_R0_addr;
  wire  mem_165_7_R0_clk;
  wire [7:0] mem_165_7_R0_data;
  wire  mem_165_7_R0_en;
  wire [25:0] mem_165_7_W0_addr;
  wire  mem_165_7_W0_clk;
  wire [7:0] mem_165_7_W0_data;
  wire  mem_165_7_W0_en;
  wire  mem_165_7_W0_mask;
  wire [25:0] mem_166_0_R0_addr;
  wire  mem_166_0_R0_clk;
  wire [7:0] mem_166_0_R0_data;
  wire  mem_166_0_R0_en;
  wire [25:0] mem_166_0_W0_addr;
  wire  mem_166_0_W0_clk;
  wire [7:0] mem_166_0_W0_data;
  wire  mem_166_0_W0_en;
  wire  mem_166_0_W0_mask;
  wire [25:0] mem_166_1_R0_addr;
  wire  mem_166_1_R0_clk;
  wire [7:0] mem_166_1_R0_data;
  wire  mem_166_1_R0_en;
  wire [25:0] mem_166_1_W0_addr;
  wire  mem_166_1_W0_clk;
  wire [7:0] mem_166_1_W0_data;
  wire  mem_166_1_W0_en;
  wire  mem_166_1_W0_mask;
  wire [25:0] mem_166_2_R0_addr;
  wire  mem_166_2_R0_clk;
  wire [7:0] mem_166_2_R0_data;
  wire  mem_166_2_R0_en;
  wire [25:0] mem_166_2_W0_addr;
  wire  mem_166_2_W0_clk;
  wire [7:0] mem_166_2_W0_data;
  wire  mem_166_2_W0_en;
  wire  mem_166_2_W0_mask;
  wire [25:0] mem_166_3_R0_addr;
  wire  mem_166_3_R0_clk;
  wire [7:0] mem_166_3_R0_data;
  wire  mem_166_3_R0_en;
  wire [25:0] mem_166_3_W0_addr;
  wire  mem_166_3_W0_clk;
  wire [7:0] mem_166_3_W0_data;
  wire  mem_166_3_W0_en;
  wire  mem_166_3_W0_mask;
  wire [25:0] mem_166_4_R0_addr;
  wire  mem_166_4_R0_clk;
  wire [7:0] mem_166_4_R0_data;
  wire  mem_166_4_R0_en;
  wire [25:0] mem_166_4_W0_addr;
  wire  mem_166_4_W0_clk;
  wire [7:0] mem_166_4_W0_data;
  wire  mem_166_4_W0_en;
  wire  mem_166_4_W0_mask;
  wire [25:0] mem_166_5_R0_addr;
  wire  mem_166_5_R0_clk;
  wire [7:0] mem_166_5_R0_data;
  wire  mem_166_5_R0_en;
  wire [25:0] mem_166_5_W0_addr;
  wire  mem_166_5_W0_clk;
  wire [7:0] mem_166_5_W0_data;
  wire  mem_166_5_W0_en;
  wire  mem_166_5_W0_mask;
  wire [25:0] mem_166_6_R0_addr;
  wire  mem_166_6_R0_clk;
  wire [7:0] mem_166_6_R0_data;
  wire  mem_166_6_R0_en;
  wire [25:0] mem_166_6_W0_addr;
  wire  mem_166_6_W0_clk;
  wire [7:0] mem_166_6_W0_data;
  wire  mem_166_6_W0_en;
  wire  mem_166_6_W0_mask;
  wire [25:0] mem_166_7_R0_addr;
  wire  mem_166_7_R0_clk;
  wire [7:0] mem_166_7_R0_data;
  wire  mem_166_7_R0_en;
  wire [25:0] mem_166_7_W0_addr;
  wire  mem_166_7_W0_clk;
  wire [7:0] mem_166_7_W0_data;
  wire  mem_166_7_W0_en;
  wire  mem_166_7_W0_mask;
  wire [25:0] mem_167_0_R0_addr;
  wire  mem_167_0_R0_clk;
  wire [7:0] mem_167_0_R0_data;
  wire  mem_167_0_R0_en;
  wire [25:0] mem_167_0_W0_addr;
  wire  mem_167_0_W0_clk;
  wire [7:0] mem_167_0_W0_data;
  wire  mem_167_0_W0_en;
  wire  mem_167_0_W0_mask;
  wire [25:0] mem_167_1_R0_addr;
  wire  mem_167_1_R0_clk;
  wire [7:0] mem_167_1_R0_data;
  wire  mem_167_1_R0_en;
  wire [25:0] mem_167_1_W0_addr;
  wire  mem_167_1_W0_clk;
  wire [7:0] mem_167_1_W0_data;
  wire  mem_167_1_W0_en;
  wire  mem_167_1_W0_mask;
  wire [25:0] mem_167_2_R0_addr;
  wire  mem_167_2_R0_clk;
  wire [7:0] mem_167_2_R0_data;
  wire  mem_167_2_R0_en;
  wire [25:0] mem_167_2_W0_addr;
  wire  mem_167_2_W0_clk;
  wire [7:0] mem_167_2_W0_data;
  wire  mem_167_2_W0_en;
  wire  mem_167_2_W0_mask;
  wire [25:0] mem_167_3_R0_addr;
  wire  mem_167_3_R0_clk;
  wire [7:0] mem_167_3_R0_data;
  wire  mem_167_3_R0_en;
  wire [25:0] mem_167_3_W0_addr;
  wire  mem_167_3_W0_clk;
  wire [7:0] mem_167_3_W0_data;
  wire  mem_167_3_W0_en;
  wire  mem_167_3_W0_mask;
  wire [25:0] mem_167_4_R0_addr;
  wire  mem_167_4_R0_clk;
  wire [7:0] mem_167_4_R0_data;
  wire  mem_167_4_R0_en;
  wire [25:0] mem_167_4_W0_addr;
  wire  mem_167_4_W0_clk;
  wire [7:0] mem_167_4_W0_data;
  wire  mem_167_4_W0_en;
  wire  mem_167_4_W0_mask;
  wire [25:0] mem_167_5_R0_addr;
  wire  mem_167_5_R0_clk;
  wire [7:0] mem_167_5_R0_data;
  wire  mem_167_5_R0_en;
  wire [25:0] mem_167_5_W0_addr;
  wire  mem_167_5_W0_clk;
  wire [7:0] mem_167_5_W0_data;
  wire  mem_167_5_W0_en;
  wire  mem_167_5_W0_mask;
  wire [25:0] mem_167_6_R0_addr;
  wire  mem_167_6_R0_clk;
  wire [7:0] mem_167_6_R0_data;
  wire  mem_167_6_R0_en;
  wire [25:0] mem_167_6_W0_addr;
  wire  mem_167_6_W0_clk;
  wire [7:0] mem_167_6_W0_data;
  wire  mem_167_6_W0_en;
  wire  mem_167_6_W0_mask;
  wire [25:0] mem_167_7_R0_addr;
  wire  mem_167_7_R0_clk;
  wire [7:0] mem_167_7_R0_data;
  wire  mem_167_7_R0_en;
  wire [25:0] mem_167_7_W0_addr;
  wire  mem_167_7_W0_clk;
  wire [7:0] mem_167_7_W0_data;
  wire  mem_167_7_W0_en;
  wire  mem_167_7_W0_mask;
  wire [25:0] mem_168_0_R0_addr;
  wire  mem_168_0_R0_clk;
  wire [7:0] mem_168_0_R0_data;
  wire  mem_168_0_R0_en;
  wire [25:0] mem_168_0_W0_addr;
  wire  mem_168_0_W0_clk;
  wire [7:0] mem_168_0_W0_data;
  wire  mem_168_0_W0_en;
  wire  mem_168_0_W0_mask;
  wire [25:0] mem_168_1_R0_addr;
  wire  mem_168_1_R0_clk;
  wire [7:0] mem_168_1_R0_data;
  wire  mem_168_1_R0_en;
  wire [25:0] mem_168_1_W0_addr;
  wire  mem_168_1_W0_clk;
  wire [7:0] mem_168_1_W0_data;
  wire  mem_168_1_W0_en;
  wire  mem_168_1_W0_mask;
  wire [25:0] mem_168_2_R0_addr;
  wire  mem_168_2_R0_clk;
  wire [7:0] mem_168_2_R0_data;
  wire  mem_168_2_R0_en;
  wire [25:0] mem_168_2_W0_addr;
  wire  mem_168_2_W0_clk;
  wire [7:0] mem_168_2_W0_data;
  wire  mem_168_2_W0_en;
  wire  mem_168_2_W0_mask;
  wire [25:0] mem_168_3_R0_addr;
  wire  mem_168_3_R0_clk;
  wire [7:0] mem_168_3_R0_data;
  wire  mem_168_3_R0_en;
  wire [25:0] mem_168_3_W0_addr;
  wire  mem_168_3_W0_clk;
  wire [7:0] mem_168_3_W0_data;
  wire  mem_168_3_W0_en;
  wire  mem_168_3_W0_mask;
  wire [25:0] mem_168_4_R0_addr;
  wire  mem_168_4_R0_clk;
  wire [7:0] mem_168_4_R0_data;
  wire  mem_168_4_R0_en;
  wire [25:0] mem_168_4_W0_addr;
  wire  mem_168_4_W0_clk;
  wire [7:0] mem_168_4_W0_data;
  wire  mem_168_4_W0_en;
  wire  mem_168_4_W0_mask;
  wire [25:0] mem_168_5_R0_addr;
  wire  mem_168_5_R0_clk;
  wire [7:0] mem_168_5_R0_data;
  wire  mem_168_5_R0_en;
  wire [25:0] mem_168_5_W0_addr;
  wire  mem_168_5_W0_clk;
  wire [7:0] mem_168_5_W0_data;
  wire  mem_168_5_W0_en;
  wire  mem_168_5_W0_mask;
  wire [25:0] mem_168_6_R0_addr;
  wire  mem_168_6_R0_clk;
  wire [7:0] mem_168_6_R0_data;
  wire  mem_168_6_R0_en;
  wire [25:0] mem_168_6_W0_addr;
  wire  mem_168_6_W0_clk;
  wire [7:0] mem_168_6_W0_data;
  wire  mem_168_6_W0_en;
  wire  mem_168_6_W0_mask;
  wire [25:0] mem_168_7_R0_addr;
  wire  mem_168_7_R0_clk;
  wire [7:0] mem_168_7_R0_data;
  wire  mem_168_7_R0_en;
  wire [25:0] mem_168_7_W0_addr;
  wire  mem_168_7_W0_clk;
  wire [7:0] mem_168_7_W0_data;
  wire  mem_168_7_W0_en;
  wire  mem_168_7_W0_mask;
  wire [25:0] mem_169_0_R0_addr;
  wire  mem_169_0_R0_clk;
  wire [7:0] mem_169_0_R0_data;
  wire  mem_169_0_R0_en;
  wire [25:0] mem_169_0_W0_addr;
  wire  mem_169_0_W0_clk;
  wire [7:0] mem_169_0_W0_data;
  wire  mem_169_0_W0_en;
  wire  mem_169_0_W0_mask;
  wire [25:0] mem_169_1_R0_addr;
  wire  mem_169_1_R0_clk;
  wire [7:0] mem_169_1_R0_data;
  wire  mem_169_1_R0_en;
  wire [25:0] mem_169_1_W0_addr;
  wire  mem_169_1_W0_clk;
  wire [7:0] mem_169_1_W0_data;
  wire  mem_169_1_W0_en;
  wire  mem_169_1_W0_mask;
  wire [25:0] mem_169_2_R0_addr;
  wire  mem_169_2_R0_clk;
  wire [7:0] mem_169_2_R0_data;
  wire  mem_169_2_R0_en;
  wire [25:0] mem_169_2_W0_addr;
  wire  mem_169_2_W0_clk;
  wire [7:0] mem_169_2_W0_data;
  wire  mem_169_2_W0_en;
  wire  mem_169_2_W0_mask;
  wire [25:0] mem_169_3_R0_addr;
  wire  mem_169_3_R0_clk;
  wire [7:0] mem_169_3_R0_data;
  wire  mem_169_3_R0_en;
  wire [25:0] mem_169_3_W0_addr;
  wire  mem_169_3_W0_clk;
  wire [7:0] mem_169_3_W0_data;
  wire  mem_169_3_W0_en;
  wire  mem_169_3_W0_mask;
  wire [25:0] mem_169_4_R0_addr;
  wire  mem_169_4_R0_clk;
  wire [7:0] mem_169_4_R0_data;
  wire  mem_169_4_R0_en;
  wire [25:0] mem_169_4_W0_addr;
  wire  mem_169_4_W0_clk;
  wire [7:0] mem_169_4_W0_data;
  wire  mem_169_4_W0_en;
  wire  mem_169_4_W0_mask;
  wire [25:0] mem_169_5_R0_addr;
  wire  mem_169_5_R0_clk;
  wire [7:0] mem_169_5_R0_data;
  wire  mem_169_5_R0_en;
  wire [25:0] mem_169_5_W0_addr;
  wire  mem_169_5_W0_clk;
  wire [7:0] mem_169_5_W0_data;
  wire  mem_169_5_W0_en;
  wire  mem_169_5_W0_mask;
  wire [25:0] mem_169_6_R0_addr;
  wire  mem_169_6_R0_clk;
  wire [7:0] mem_169_6_R0_data;
  wire  mem_169_6_R0_en;
  wire [25:0] mem_169_6_W0_addr;
  wire  mem_169_6_W0_clk;
  wire [7:0] mem_169_6_W0_data;
  wire  mem_169_6_W0_en;
  wire  mem_169_6_W0_mask;
  wire [25:0] mem_169_7_R0_addr;
  wire  mem_169_7_R0_clk;
  wire [7:0] mem_169_7_R0_data;
  wire  mem_169_7_R0_en;
  wire [25:0] mem_169_7_W0_addr;
  wire  mem_169_7_W0_clk;
  wire [7:0] mem_169_7_W0_data;
  wire  mem_169_7_W0_en;
  wire  mem_169_7_W0_mask;
  wire [25:0] mem_170_0_R0_addr;
  wire  mem_170_0_R0_clk;
  wire [7:0] mem_170_0_R0_data;
  wire  mem_170_0_R0_en;
  wire [25:0] mem_170_0_W0_addr;
  wire  mem_170_0_W0_clk;
  wire [7:0] mem_170_0_W0_data;
  wire  mem_170_0_W0_en;
  wire  mem_170_0_W0_mask;
  wire [25:0] mem_170_1_R0_addr;
  wire  mem_170_1_R0_clk;
  wire [7:0] mem_170_1_R0_data;
  wire  mem_170_1_R0_en;
  wire [25:0] mem_170_1_W0_addr;
  wire  mem_170_1_W0_clk;
  wire [7:0] mem_170_1_W0_data;
  wire  mem_170_1_W0_en;
  wire  mem_170_1_W0_mask;
  wire [25:0] mem_170_2_R0_addr;
  wire  mem_170_2_R0_clk;
  wire [7:0] mem_170_2_R0_data;
  wire  mem_170_2_R0_en;
  wire [25:0] mem_170_2_W0_addr;
  wire  mem_170_2_W0_clk;
  wire [7:0] mem_170_2_W0_data;
  wire  mem_170_2_W0_en;
  wire  mem_170_2_W0_mask;
  wire [25:0] mem_170_3_R0_addr;
  wire  mem_170_3_R0_clk;
  wire [7:0] mem_170_3_R0_data;
  wire  mem_170_3_R0_en;
  wire [25:0] mem_170_3_W0_addr;
  wire  mem_170_3_W0_clk;
  wire [7:0] mem_170_3_W0_data;
  wire  mem_170_3_W0_en;
  wire  mem_170_3_W0_mask;
  wire [25:0] mem_170_4_R0_addr;
  wire  mem_170_4_R0_clk;
  wire [7:0] mem_170_4_R0_data;
  wire  mem_170_4_R0_en;
  wire [25:0] mem_170_4_W0_addr;
  wire  mem_170_4_W0_clk;
  wire [7:0] mem_170_4_W0_data;
  wire  mem_170_4_W0_en;
  wire  mem_170_4_W0_mask;
  wire [25:0] mem_170_5_R0_addr;
  wire  mem_170_5_R0_clk;
  wire [7:0] mem_170_5_R0_data;
  wire  mem_170_5_R0_en;
  wire [25:0] mem_170_5_W0_addr;
  wire  mem_170_5_W0_clk;
  wire [7:0] mem_170_5_W0_data;
  wire  mem_170_5_W0_en;
  wire  mem_170_5_W0_mask;
  wire [25:0] mem_170_6_R0_addr;
  wire  mem_170_6_R0_clk;
  wire [7:0] mem_170_6_R0_data;
  wire  mem_170_6_R0_en;
  wire [25:0] mem_170_6_W0_addr;
  wire  mem_170_6_W0_clk;
  wire [7:0] mem_170_6_W0_data;
  wire  mem_170_6_W0_en;
  wire  mem_170_6_W0_mask;
  wire [25:0] mem_170_7_R0_addr;
  wire  mem_170_7_R0_clk;
  wire [7:0] mem_170_7_R0_data;
  wire  mem_170_7_R0_en;
  wire [25:0] mem_170_7_W0_addr;
  wire  mem_170_7_W0_clk;
  wire [7:0] mem_170_7_W0_data;
  wire  mem_170_7_W0_en;
  wire  mem_170_7_W0_mask;
  wire [25:0] mem_171_0_R0_addr;
  wire  mem_171_0_R0_clk;
  wire [7:0] mem_171_0_R0_data;
  wire  mem_171_0_R0_en;
  wire [25:0] mem_171_0_W0_addr;
  wire  mem_171_0_W0_clk;
  wire [7:0] mem_171_0_W0_data;
  wire  mem_171_0_W0_en;
  wire  mem_171_0_W0_mask;
  wire [25:0] mem_171_1_R0_addr;
  wire  mem_171_1_R0_clk;
  wire [7:0] mem_171_1_R0_data;
  wire  mem_171_1_R0_en;
  wire [25:0] mem_171_1_W0_addr;
  wire  mem_171_1_W0_clk;
  wire [7:0] mem_171_1_W0_data;
  wire  mem_171_1_W0_en;
  wire  mem_171_1_W0_mask;
  wire [25:0] mem_171_2_R0_addr;
  wire  mem_171_2_R0_clk;
  wire [7:0] mem_171_2_R0_data;
  wire  mem_171_2_R0_en;
  wire [25:0] mem_171_2_W0_addr;
  wire  mem_171_2_W0_clk;
  wire [7:0] mem_171_2_W0_data;
  wire  mem_171_2_W0_en;
  wire  mem_171_2_W0_mask;
  wire [25:0] mem_171_3_R0_addr;
  wire  mem_171_3_R0_clk;
  wire [7:0] mem_171_3_R0_data;
  wire  mem_171_3_R0_en;
  wire [25:0] mem_171_3_W0_addr;
  wire  mem_171_3_W0_clk;
  wire [7:0] mem_171_3_W0_data;
  wire  mem_171_3_W0_en;
  wire  mem_171_3_W0_mask;
  wire [25:0] mem_171_4_R0_addr;
  wire  mem_171_4_R0_clk;
  wire [7:0] mem_171_4_R0_data;
  wire  mem_171_4_R0_en;
  wire [25:0] mem_171_4_W0_addr;
  wire  mem_171_4_W0_clk;
  wire [7:0] mem_171_4_W0_data;
  wire  mem_171_4_W0_en;
  wire  mem_171_4_W0_mask;
  wire [25:0] mem_171_5_R0_addr;
  wire  mem_171_5_R0_clk;
  wire [7:0] mem_171_5_R0_data;
  wire  mem_171_5_R0_en;
  wire [25:0] mem_171_5_W0_addr;
  wire  mem_171_5_W0_clk;
  wire [7:0] mem_171_5_W0_data;
  wire  mem_171_5_W0_en;
  wire  mem_171_5_W0_mask;
  wire [25:0] mem_171_6_R0_addr;
  wire  mem_171_6_R0_clk;
  wire [7:0] mem_171_6_R0_data;
  wire  mem_171_6_R0_en;
  wire [25:0] mem_171_6_W0_addr;
  wire  mem_171_6_W0_clk;
  wire [7:0] mem_171_6_W0_data;
  wire  mem_171_6_W0_en;
  wire  mem_171_6_W0_mask;
  wire [25:0] mem_171_7_R0_addr;
  wire  mem_171_7_R0_clk;
  wire [7:0] mem_171_7_R0_data;
  wire  mem_171_7_R0_en;
  wire [25:0] mem_171_7_W0_addr;
  wire  mem_171_7_W0_clk;
  wire [7:0] mem_171_7_W0_data;
  wire  mem_171_7_W0_en;
  wire  mem_171_7_W0_mask;
  wire [25:0] mem_172_0_R0_addr;
  wire  mem_172_0_R0_clk;
  wire [7:0] mem_172_0_R0_data;
  wire  mem_172_0_R0_en;
  wire [25:0] mem_172_0_W0_addr;
  wire  mem_172_0_W0_clk;
  wire [7:0] mem_172_0_W0_data;
  wire  mem_172_0_W0_en;
  wire  mem_172_0_W0_mask;
  wire [25:0] mem_172_1_R0_addr;
  wire  mem_172_1_R0_clk;
  wire [7:0] mem_172_1_R0_data;
  wire  mem_172_1_R0_en;
  wire [25:0] mem_172_1_W0_addr;
  wire  mem_172_1_W0_clk;
  wire [7:0] mem_172_1_W0_data;
  wire  mem_172_1_W0_en;
  wire  mem_172_1_W0_mask;
  wire [25:0] mem_172_2_R0_addr;
  wire  mem_172_2_R0_clk;
  wire [7:0] mem_172_2_R0_data;
  wire  mem_172_2_R0_en;
  wire [25:0] mem_172_2_W0_addr;
  wire  mem_172_2_W0_clk;
  wire [7:0] mem_172_2_W0_data;
  wire  mem_172_2_W0_en;
  wire  mem_172_2_W0_mask;
  wire [25:0] mem_172_3_R0_addr;
  wire  mem_172_3_R0_clk;
  wire [7:0] mem_172_3_R0_data;
  wire  mem_172_3_R0_en;
  wire [25:0] mem_172_3_W0_addr;
  wire  mem_172_3_W0_clk;
  wire [7:0] mem_172_3_W0_data;
  wire  mem_172_3_W0_en;
  wire  mem_172_3_W0_mask;
  wire [25:0] mem_172_4_R0_addr;
  wire  mem_172_4_R0_clk;
  wire [7:0] mem_172_4_R0_data;
  wire  mem_172_4_R0_en;
  wire [25:0] mem_172_4_W0_addr;
  wire  mem_172_4_W0_clk;
  wire [7:0] mem_172_4_W0_data;
  wire  mem_172_4_W0_en;
  wire  mem_172_4_W0_mask;
  wire [25:0] mem_172_5_R0_addr;
  wire  mem_172_5_R0_clk;
  wire [7:0] mem_172_5_R0_data;
  wire  mem_172_5_R0_en;
  wire [25:0] mem_172_5_W0_addr;
  wire  mem_172_5_W0_clk;
  wire [7:0] mem_172_5_W0_data;
  wire  mem_172_5_W0_en;
  wire  mem_172_5_W0_mask;
  wire [25:0] mem_172_6_R0_addr;
  wire  mem_172_6_R0_clk;
  wire [7:0] mem_172_6_R0_data;
  wire  mem_172_6_R0_en;
  wire [25:0] mem_172_6_W0_addr;
  wire  mem_172_6_W0_clk;
  wire [7:0] mem_172_6_W0_data;
  wire  mem_172_6_W0_en;
  wire  mem_172_6_W0_mask;
  wire [25:0] mem_172_7_R0_addr;
  wire  mem_172_7_R0_clk;
  wire [7:0] mem_172_7_R0_data;
  wire  mem_172_7_R0_en;
  wire [25:0] mem_172_7_W0_addr;
  wire  mem_172_7_W0_clk;
  wire [7:0] mem_172_7_W0_data;
  wire  mem_172_7_W0_en;
  wire  mem_172_7_W0_mask;
  wire [25:0] mem_173_0_R0_addr;
  wire  mem_173_0_R0_clk;
  wire [7:0] mem_173_0_R0_data;
  wire  mem_173_0_R0_en;
  wire [25:0] mem_173_0_W0_addr;
  wire  mem_173_0_W0_clk;
  wire [7:0] mem_173_0_W0_data;
  wire  mem_173_0_W0_en;
  wire  mem_173_0_W0_mask;
  wire [25:0] mem_173_1_R0_addr;
  wire  mem_173_1_R0_clk;
  wire [7:0] mem_173_1_R0_data;
  wire  mem_173_1_R0_en;
  wire [25:0] mem_173_1_W0_addr;
  wire  mem_173_1_W0_clk;
  wire [7:0] mem_173_1_W0_data;
  wire  mem_173_1_W0_en;
  wire  mem_173_1_W0_mask;
  wire [25:0] mem_173_2_R0_addr;
  wire  mem_173_2_R0_clk;
  wire [7:0] mem_173_2_R0_data;
  wire  mem_173_2_R0_en;
  wire [25:0] mem_173_2_W0_addr;
  wire  mem_173_2_W0_clk;
  wire [7:0] mem_173_2_W0_data;
  wire  mem_173_2_W0_en;
  wire  mem_173_2_W0_mask;
  wire [25:0] mem_173_3_R0_addr;
  wire  mem_173_3_R0_clk;
  wire [7:0] mem_173_3_R0_data;
  wire  mem_173_3_R0_en;
  wire [25:0] mem_173_3_W0_addr;
  wire  mem_173_3_W0_clk;
  wire [7:0] mem_173_3_W0_data;
  wire  mem_173_3_W0_en;
  wire  mem_173_3_W0_mask;
  wire [25:0] mem_173_4_R0_addr;
  wire  mem_173_4_R0_clk;
  wire [7:0] mem_173_4_R0_data;
  wire  mem_173_4_R0_en;
  wire [25:0] mem_173_4_W0_addr;
  wire  mem_173_4_W0_clk;
  wire [7:0] mem_173_4_W0_data;
  wire  mem_173_4_W0_en;
  wire  mem_173_4_W0_mask;
  wire [25:0] mem_173_5_R0_addr;
  wire  mem_173_5_R0_clk;
  wire [7:0] mem_173_5_R0_data;
  wire  mem_173_5_R0_en;
  wire [25:0] mem_173_5_W0_addr;
  wire  mem_173_5_W0_clk;
  wire [7:0] mem_173_5_W0_data;
  wire  mem_173_5_W0_en;
  wire  mem_173_5_W0_mask;
  wire [25:0] mem_173_6_R0_addr;
  wire  mem_173_6_R0_clk;
  wire [7:0] mem_173_6_R0_data;
  wire  mem_173_6_R0_en;
  wire [25:0] mem_173_6_W0_addr;
  wire  mem_173_6_W0_clk;
  wire [7:0] mem_173_6_W0_data;
  wire  mem_173_6_W0_en;
  wire  mem_173_6_W0_mask;
  wire [25:0] mem_173_7_R0_addr;
  wire  mem_173_7_R0_clk;
  wire [7:0] mem_173_7_R0_data;
  wire  mem_173_7_R0_en;
  wire [25:0] mem_173_7_W0_addr;
  wire  mem_173_7_W0_clk;
  wire [7:0] mem_173_7_W0_data;
  wire  mem_173_7_W0_en;
  wire  mem_173_7_W0_mask;
  wire [25:0] mem_174_0_R0_addr;
  wire  mem_174_0_R0_clk;
  wire [7:0] mem_174_0_R0_data;
  wire  mem_174_0_R0_en;
  wire [25:0] mem_174_0_W0_addr;
  wire  mem_174_0_W0_clk;
  wire [7:0] mem_174_0_W0_data;
  wire  mem_174_0_W0_en;
  wire  mem_174_0_W0_mask;
  wire [25:0] mem_174_1_R0_addr;
  wire  mem_174_1_R0_clk;
  wire [7:0] mem_174_1_R0_data;
  wire  mem_174_1_R0_en;
  wire [25:0] mem_174_1_W0_addr;
  wire  mem_174_1_W0_clk;
  wire [7:0] mem_174_1_W0_data;
  wire  mem_174_1_W0_en;
  wire  mem_174_1_W0_mask;
  wire [25:0] mem_174_2_R0_addr;
  wire  mem_174_2_R0_clk;
  wire [7:0] mem_174_2_R0_data;
  wire  mem_174_2_R0_en;
  wire [25:0] mem_174_2_W0_addr;
  wire  mem_174_2_W0_clk;
  wire [7:0] mem_174_2_W0_data;
  wire  mem_174_2_W0_en;
  wire  mem_174_2_W0_mask;
  wire [25:0] mem_174_3_R0_addr;
  wire  mem_174_3_R0_clk;
  wire [7:0] mem_174_3_R0_data;
  wire  mem_174_3_R0_en;
  wire [25:0] mem_174_3_W0_addr;
  wire  mem_174_3_W0_clk;
  wire [7:0] mem_174_3_W0_data;
  wire  mem_174_3_W0_en;
  wire  mem_174_3_W0_mask;
  wire [25:0] mem_174_4_R0_addr;
  wire  mem_174_4_R0_clk;
  wire [7:0] mem_174_4_R0_data;
  wire  mem_174_4_R0_en;
  wire [25:0] mem_174_4_W0_addr;
  wire  mem_174_4_W0_clk;
  wire [7:0] mem_174_4_W0_data;
  wire  mem_174_4_W0_en;
  wire  mem_174_4_W0_mask;
  wire [25:0] mem_174_5_R0_addr;
  wire  mem_174_5_R0_clk;
  wire [7:0] mem_174_5_R0_data;
  wire  mem_174_5_R0_en;
  wire [25:0] mem_174_5_W0_addr;
  wire  mem_174_5_W0_clk;
  wire [7:0] mem_174_5_W0_data;
  wire  mem_174_5_W0_en;
  wire  mem_174_5_W0_mask;
  wire [25:0] mem_174_6_R0_addr;
  wire  mem_174_6_R0_clk;
  wire [7:0] mem_174_6_R0_data;
  wire  mem_174_6_R0_en;
  wire [25:0] mem_174_6_W0_addr;
  wire  mem_174_6_W0_clk;
  wire [7:0] mem_174_6_W0_data;
  wire  mem_174_6_W0_en;
  wire  mem_174_6_W0_mask;
  wire [25:0] mem_174_7_R0_addr;
  wire  mem_174_7_R0_clk;
  wire [7:0] mem_174_7_R0_data;
  wire  mem_174_7_R0_en;
  wire [25:0] mem_174_7_W0_addr;
  wire  mem_174_7_W0_clk;
  wire [7:0] mem_174_7_W0_data;
  wire  mem_174_7_W0_en;
  wire  mem_174_7_W0_mask;
  wire [25:0] mem_175_0_R0_addr;
  wire  mem_175_0_R0_clk;
  wire [7:0] mem_175_0_R0_data;
  wire  mem_175_0_R0_en;
  wire [25:0] mem_175_0_W0_addr;
  wire  mem_175_0_W0_clk;
  wire [7:0] mem_175_0_W0_data;
  wire  mem_175_0_W0_en;
  wire  mem_175_0_W0_mask;
  wire [25:0] mem_175_1_R0_addr;
  wire  mem_175_1_R0_clk;
  wire [7:0] mem_175_1_R0_data;
  wire  mem_175_1_R0_en;
  wire [25:0] mem_175_1_W0_addr;
  wire  mem_175_1_W0_clk;
  wire [7:0] mem_175_1_W0_data;
  wire  mem_175_1_W0_en;
  wire  mem_175_1_W0_mask;
  wire [25:0] mem_175_2_R0_addr;
  wire  mem_175_2_R0_clk;
  wire [7:0] mem_175_2_R0_data;
  wire  mem_175_2_R0_en;
  wire [25:0] mem_175_2_W0_addr;
  wire  mem_175_2_W0_clk;
  wire [7:0] mem_175_2_W0_data;
  wire  mem_175_2_W0_en;
  wire  mem_175_2_W0_mask;
  wire [25:0] mem_175_3_R0_addr;
  wire  mem_175_3_R0_clk;
  wire [7:0] mem_175_3_R0_data;
  wire  mem_175_3_R0_en;
  wire [25:0] mem_175_3_W0_addr;
  wire  mem_175_3_W0_clk;
  wire [7:0] mem_175_3_W0_data;
  wire  mem_175_3_W0_en;
  wire  mem_175_3_W0_mask;
  wire [25:0] mem_175_4_R0_addr;
  wire  mem_175_4_R0_clk;
  wire [7:0] mem_175_4_R0_data;
  wire  mem_175_4_R0_en;
  wire [25:0] mem_175_4_W0_addr;
  wire  mem_175_4_W0_clk;
  wire [7:0] mem_175_4_W0_data;
  wire  mem_175_4_W0_en;
  wire  mem_175_4_W0_mask;
  wire [25:0] mem_175_5_R0_addr;
  wire  mem_175_5_R0_clk;
  wire [7:0] mem_175_5_R0_data;
  wire  mem_175_5_R0_en;
  wire [25:0] mem_175_5_W0_addr;
  wire  mem_175_5_W0_clk;
  wire [7:0] mem_175_5_W0_data;
  wire  mem_175_5_W0_en;
  wire  mem_175_5_W0_mask;
  wire [25:0] mem_175_6_R0_addr;
  wire  mem_175_6_R0_clk;
  wire [7:0] mem_175_6_R0_data;
  wire  mem_175_6_R0_en;
  wire [25:0] mem_175_6_W0_addr;
  wire  mem_175_6_W0_clk;
  wire [7:0] mem_175_6_W0_data;
  wire  mem_175_6_W0_en;
  wire  mem_175_6_W0_mask;
  wire [25:0] mem_175_7_R0_addr;
  wire  mem_175_7_R0_clk;
  wire [7:0] mem_175_7_R0_data;
  wire  mem_175_7_R0_en;
  wire [25:0] mem_175_7_W0_addr;
  wire  mem_175_7_W0_clk;
  wire [7:0] mem_175_7_W0_data;
  wire  mem_175_7_W0_en;
  wire  mem_175_7_W0_mask;
  wire [25:0] mem_176_0_R0_addr;
  wire  mem_176_0_R0_clk;
  wire [7:0] mem_176_0_R0_data;
  wire  mem_176_0_R0_en;
  wire [25:0] mem_176_0_W0_addr;
  wire  mem_176_0_W0_clk;
  wire [7:0] mem_176_0_W0_data;
  wire  mem_176_0_W0_en;
  wire  mem_176_0_W0_mask;
  wire [25:0] mem_176_1_R0_addr;
  wire  mem_176_1_R0_clk;
  wire [7:0] mem_176_1_R0_data;
  wire  mem_176_1_R0_en;
  wire [25:0] mem_176_1_W0_addr;
  wire  mem_176_1_W0_clk;
  wire [7:0] mem_176_1_W0_data;
  wire  mem_176_1_W0_en;
  wire  mem_176_1_W0_mask;
  wire [25:0] mem_176_2_R0_addr;
  wire  mem_176_2_R0_clk;
  wire [7:0] mem_176_2_R0_data;
  wire  mem_176_2_R0_en;
  wire [25:0] mem_176_2_W0_addr;
  wire  mem_176_2_W0_clk;
  wire [7:0] mem_176_2_W0_data;
  wire  mem_176_2_W0_en;
  wire  mem_176_2_W0_mask;
  wire [25:0] mem_176_3_R0_addr;
  wire  mem_176_3_R0_clk;
  wire [7:0] mem_176_3_R0_data;
  wire  mem_176_3_R0_en;
  wire [25:0] mem_176_3_W0_addr;
  wire  mem_176_3_W0_clk;
  wire [7:0] mem_176_3_W0_data;
  wire  mem_176_3_W0_en;
  wire  mem_176_3_W0_mask;
  wire [25:0] mem_176_4_R0_addr;
  wire  mem_176_4_R0_clk;
  wire [7:0] mem_176_4_R0_data;
  wire  mem_176_4_R0_en;
  wire [25:0] mem_176_4_W0_addr;
  wire  mem_176_4_W0_clk;
  wire [7:0] mem_176_4_W0_data;
  wire  mem_176_4_W0_en;
  wire  mem_176_4_W0_mask;
  wire [25:0] mem_176_5_R0_addr;
  wire  mem_176_5_R0_clk;
  wire [7:0] mem_176_5_R0_data;
  wire  mem_176_5_R0_en;
  wire [25:0] mem_176_5_W0_addr;
  wire  mem_176_5_W0_clk;
  wire [7:0] mem_176_5_W0_data;
  wire  mem_176_5_W0_en;
  wire  mem_176_5_W0_mask;
  wire [25:0] mem_176_6_R0_addr;
  wire  mem_176_6_R0_clk;
  wire [7:0] mem_176_6_R0_data;
  wire  mem_176_6_R0_en;
  wire [25:0] mem_176_6_W0_addr;
  wire  mem_176_6_W0_clk;
  wire [7:0] mem_176_6_W0_data;
  wire  mem_176_6_W0_en;
  wire  mem_176_6_W0_mask;
  wire [25:0] mem_176_7_R0_addr;
  wire  mem_176_7_R0_clk;
  wire [7:0] mem_176_7_R0_data;
  wire  mem_176_7_R0_en;
  wire [25:0] mem_176_7_W0_addr;
  wire  mem_176_7_W0_clk;
  wire [7:0] mem_176_7_W0_data;
  wire  mem_176_7_W0_en;
  wire  mem_176_7_W0_mask;
  wire [25:0] mem_177_0_R0_addr;
  wire  mem_177_0_R0_clk;
  wire [7:0] mem_177_0_R0_data;
  wire  mem_177_0_R0_en;
  wire [25:0] mem_177_0_W0_addr;
  wire  mem_177_0_W0_clk;
  wire [7:0] mem_177_0_W0_data;
  wire  mem_177_0_W0_en;
  wire  mem_177_0_W0_mask;
  wire [25:0] mem_177_1_R0_addr;
  wire  mem_177_1_R0_clk;
  wire [7:0] mem_177_1_R0_data;
  wire  mem_177_1_R0_en;
  wire [25:0] mem_177_1_W0_addr;
  wire  mem_177_1_W0_clk;
  wire [7:0] mem_177_1_W0_data;
  wire  mem_177_1_W0_en;
  wire  mem_177_1_W0_mask;
  wire [25:0] mem_177_2_R0_addr;
  wire  mem_177_2_R0_clk;
  wire [7:0] mem_177_2_R0_data;
  wire  mem_177_2_R0_en;
  wire [25:0] mem_177_2_W0_addr;
  wire  mem_177_2_W0_clk;
  wire [7:0] mem_177_2_W0_data;
  wire  mem_177_2_W0_en;
  wire  mem_177_2_W0_mask;
  wire [25:0] mem_177_3_R0_addr;
  wire  mem_177_3_R0_clk;
  wire [7:0] mem_177_3_R0_data;
  wire  mem_177_3_R0_en;
  wire [25:0] mem_177_3_W0_addr;
  wire  mem_177_3_W0_clk;
  wire [7:0] mem_177_3_W0_data;
  wire  mem_177_3_W0_en;
  wire  mem_177_3_W0_mask;
  wire [25:0] mem_177_4_R0_addr;
  wire  mem_177_4_R0_clk;
  wire [7:0] mem_177_4_R0_data;
  wire  mem_177_4_R0_en;
  wire [25:0] mem_177_4_W0_addr;
  wire  mem_177_4_W0_clk;
  wire [7:0] mem_177_4_W0_data;
  wire  mem_177_4_W0_en;
  wire  mem_177_4_W0_mask;
  wire [25:0] mem_177_5_R0_addr;
  wire  mem_177_5_R0_clk;
  wire [7:0] mem_177_5_R0_data;
  wire  mem_177_5_R0_en;
  wire [25:0] mem_177_5_W0_addr;
  wire  mem_177_5_W0_clk;
  wire [7:0] mem_177_5_W0_data;
  wire  mem_177_5_W0_en;
  wire  mem_177_5_W0_mask;
  wire [25:0] mem_177_6_R0_addr;
  wire  mem_177_6_R0_clk;
  wire [7:0] mem_177_6_R0_data;
  wire  mem_177_6_R0_en;
  wire [25:0] mem_177_6_W0_addr;
  wire  mem_177_6_W0_clk;
  wire [7:0] mem_177_6_W0_data;
  wire  mem_177_6_W0_en;
  wire  mem_177_6_W0_mask;
  wire [25:0] mem_177_7_R0_addr;
  wire  mem_177_7_R0_clk;
  wire [7:0] mem_177_7_R0_data;
  wire  mem_177_7_R0_en;
  wire [25:0] mem_177_7_W0_addr;
  wire  mem_177_7_W0_clk;
  wire [7:0] mem_177_7_W0_data;
  wire  mem_177_7_W0_en;
  wire  mem_177_7_W0_mask;
  wire [25:0] mem_178_0_R0_addr;
  wire  mem_178_0_R0_clk;
  wire [7:0] mem_178_0_R0_data;
  wire  mem_178_0_R0_en;
  wire [25:0] mem_178_0_W0_addr;
  wire  mem_178_0_W0_clk;
  wire [7:0] mem_178_0_W0_data;
  wire  mem_178_0_W0_en;
  wire  mem_178_0_W0_mask;
  wire [25:0] mem_178_1_R0_addr;
  wire  mem_178_1_R0_clk;
  wire [7:0] mem_178_1_R0_data;
  wire  mem_178_1_R0_en;
  wire [25:0] mem_178_1_W0_addr;
  wire  mem_178_1_W0_clk;
  wire [7:0] mem_178_1_W0_data;
  wire  mem_178_1_W0_en;
  wire  mem_178_1_W0_mask;
  wire [25:0] mem_178_2_R0_addr;
  wire  mem_178_2_R0_clk;
  wire [7:0] mem_178_2_R0_data;
  wire  mem_178_2_R0_en;
  wire [25:0] mem_178_2_W0_addr;
  wire  mem_178_2_W0_clk;
  wire [7:0] mem_178_2_W0_data;
  wire  mem_178_2_W0_en;
  wire  mem_178_2_W0_mask;
  wire [25:0] mem_178_3_R0_addr;
  wire  mem_178_3_R0_clk;
  wire [7:0] mem_178_3_R0_data;
  wire  mem_178_3_R0_en;
  wire [25:0] mem_178_3_W0_addr;
  wire  mem_178_3_W0_clk;
  wire [7:0] mem_178_3_W0_data;
  wire  mem_178_3_W0_en;
  wire  mem_178_3_W0_mask;
  wire [25:0] mem_178_4_R0_addr;
  wire  mem_178_4_R0_clk;
  wire [7:0] mem_178_4_R0_data;
  wire  mem_178_4_R0_en;
  wire [25:0] mem_178_4_W0_addr;
  wire  mem_178_4_W0_clk;
  wire [7:0] mem_178_4_W0_data;
  wire  mem_178_4_W0_en;
  wire  mem_178_4_W0_mask;
  wire [25:0] mem_178_5_R0_addr;
  wire  mem_178_5_R0_clk;
  wire [7:0] mem_178_5_R0_data;
  wire  mem_178_5_R0_en;
  wire [25:0] mem_178_5_W0_addr;
  wire  mem_178_5_W0_clk;
  wire [7:0] mem_178_5_W0_data;
  wire  mem_178_5_W0_en;
  wire  mem_178_5_W0_mask;
  wire [25:0] mem_178_6_R0_addr;
  wire  mem_178_6_R0_clk;
  wire [7:0] mem_178_6_R0_data;
  wire  mem_178_6_R0_en;
  wire [25:0] mem_178_6_W0_addr;
  wire  mem_178_6_W0_clk;
  wire [7:0] mem_178_6_W0_data;
  wire  mem_178_6_W0_en;
  wire  mem_178_6_W0_mask;
  wire [25:0] mem_178_7_R0_addr;
  wire  mem_178_7_R0_clk;
  wire [7:0] mem_178_7_R0_data;
  wire  mem_178_7_R0_en;
  wire [25:0] mem_178_7_W0_addr;
  wire  mem_178_7_W0_clk;
  wire [7:0] mem_178_7_W0_data;
  wire  mem_178_7_W0_en;
  wire  mem_178_7_W0_mask;
  wire [25:0] mem_179_0_R0_addr;
  wire  mem_179_0_R0_clk;
  wire [7:0] mem_179_0_R0_data;
  wire  mem_179_0_R0_en;
  wire [25:0] mem_179_0_W0_addr;
  wire  mem_179_0_W0_clk;
  wire [7:0] mem_179_0_W0_data;
  wire  mem_179_0_W0_en;
  wire  mem_179_0_W0_mask;
  wire [25:0] mem_179_1_R0_addr;
  wire  mem_179_1_R0_clk;
  wire [7:0] mem_179_1_R0_data;
  wire  mem_179_1_R0_en;
  wire [25:0] mem_179_1_W0_addr;
  wire  mem_179_1_W0_clk;
  wire [7:0] mem_179_1_W0_data;
  wire  mem_179_1_W0_en;
  wire  mem_179_1_W0_mask;
  wire [25:0] mem_179_2_R0_addr;
  wire  mem_179_2_R0_clk;
  wire [7:0] mem_179_2_R0_data;
  wire  mem_179_2_R0_en;
  wire [25:0] mem_179_2_W0_addr;
  wire  mem_179_2_W0_clk;
  wire [7:0] mem_179_2_W0_data;
  wire  mem_179_2_W0_en;
  wire  mem_179_2_W0_mask;
  wire [25:0] mem_179_3_R0_addr;
  wire  mem_179_3_R0_clk;
  wire [7:0] mem_179_3_R0_data;
  wire  mem_179_3_R0_en;
  wire [25:0] mem_179_3_W0_addr;
  wire  mem_179_3_W0_clk;
  wire [7:0] mem_179_3_W0_data;
  wire  mem_179_3_W0_en;
  wire  mem_179_3_W0_mask;
  wire [25:0] mem_179_4_R0_addr;
  wire  mem_179_4_R0_clk;
  wire [7:0] mem_179_4_R0_data;
  wire  mem_179_4_R0_en;
  wire [25:0] mem_179_4_W0_addr;
  wire  mem_179_4_W0_clk;
  wire [7:0] mem_179_4_W0_data;
  wire  mem_179_4_W0_en;
  wire  mem_179_4_W0_mask;
  wire [25:0] mem_179_5_R0_addr;
  wire  mem_179_5_R0_clk;
  wire [7:0] mem_179_5_R0_data;
  wire  mem_179_5_R0_en;
  wire [25:0] mem_179_5_W0_addr;
  wire  mem_179_5_W0_clk;
  wire [7:0] mem_179_5_W0_data;
  wire  mem_179_5_W0_en;
  wire  mem_179_5_W0_mask;
  wire [25:0] mem_179_6_R0_addr;
  wire  mem_179_6_R0_clk;
  wire [7:0] mem_179_6_R0_data;
  wire  mem_179_6_R0_en;
  wire [25:0] mem_179_6_W0_addr;
  wire  mem_179_6_W0_clk;
  wire [7:0] mem_179_6_W0_data;
  wire  mem_179_6_W0_en;
  wire  mem_179_6_W0_mask;
  wire [25:0] mem_179_7_R0_addr;
  wire  mem_179_7_R0_clk;
  wire [7:0] mem_179_7_R0_data;
  wire  mem_179_7_R0_en;
  wire [25:0] mem_179_7_W0_addr;
  wire  mem_179_7_W0_clk;
  wire [7:0] mem_179_7_W0_data;
  wire  mem_179_7_W0_en;
  wire  mem_179_7_W0_mask;
  wire [25:0] mem_180_0_R0_addr;
  wire  mem_180_0_R0_clk;
  wire [7:0] mem_180_0_R0_data;
  wire  mem_180_0_R0_en;
  wire [25:0] mem_180_0_W0_addr;
  wire  mem_180_0_W0_clk;
  wire [7:0] mem_180_0_W0_data;
  wire  mem_180_0_W0_en;
  wire  mem_180_0_W0_mask;
  wire [25:0] mem_180_1_R0_addr;
  wire  mem_180_1_R0_clk;
  wire [7:0] mem_180_1_R0_data;
  wire  mem_180_1_R0_en;
  wire [25:0] mem_180_1_W0_addr;
  wire  mem_180_1_W0_clk;
  wire [7:0] mem_180_1_W0_data;
  wire  mem_180_1_W0_en;
  wire  mem_180_1_W0_mask;
  wire [25:0] mem_180_2_R0_addr;
  wire  mem_180_2_R0_clk;
  wire [7:0] mem_180_2_R0_data;
  wire  mem_180_2_R0_en;
  wire [25:0] mem_180_2_W0_addr;
  wire  mem_180_2_W0_clk;
  wire [7:0] mem_180_2_W0_data;
  wire  mem_180_2_W0_en;
  wire  mem_180_2_W0_mask;
  wire [25:0] mem_180_3_R0_addr;
  wire  mem_180_3_R0_clk;
  wire [7:0] mem_180_3_R0_data;
  wire  mem_180_3_R0_en;
  wire [25:0] mem_180_3_W0_addr;
  wire  mem_180_3_W0_clk;
  wire [7:0] mem_180_3_W0_data;
  wire  mem_180_3_W0_en;
  wire  mem_180_3_W0_mask;
  wire [25:0] mem_180_4_R0_addr;
  wire  mem_180_4_R0_clk;
  wire [7:0] mem_180_4_R0_data;
  wire  mem_180_4_R0_en;
  wire [25:0] mem_180_4_W0_addr;
  wire  mem_180_4_W0_clk;
  wire [7:0] mem_180_4_W0_data;
  wire  mem_180_4_W0_en;
  wire  mem_180_4_W0_mask;
  wire [25:0] mem_180_5_R0_addr;
  wire  mem_180_5_R0_clk;
  wire [7:0] mem_180_5_R0_data;
  wire  mem_180_5_R0_en;
  wire [25:0] mem_180_5_W0_addr;
  wire  mem_180_5_W0_clk;
  wire [7:0] mem_180_5_W0_data;
  wire  mem_180_5_W0_en;
  wire  mem_180_5_W0_mask;
  wire [25:0] mem_180_6_R0_addr;
  wire  mem_180_6_R0_clk;
  wire [7:0] mem_180_6_R0_data;
  wire  mem_180_6_R0_en;
  wire [25:0] mem_180_6_W0_addr;
  wire  mem_180_6_W0_clk;
  wire [7:0] mem_180_6_W0_data;
  wire  mem_180_6_W0_en;
  wire  mem_180_6_W0_mask;
  wire [25:0] mem_180_7_R0_addr;
  wire  mem_180_7_R0_clk;
  wire [7:0] mem_180_7_R0_data;
  wire  mem_180_7_R0_en;
  wire [25:0] mem_180_7_W0_addr;
  wire  mem_180_7_W0_clk;
  wire [7:0] mem_180_7_W0_data;
  wire  mem_180_7_W0_en;
  wire  mem_180_7_W0_mask;
  wire [25:0] mem_181_0_R0_addr;
  wire  mem_181_0_R0_clk;
  wire [7:0] mem_181_0_R0_data;
  wire  mem_181_0_R0_en;
  wire [25:0] mem_181_0_W0_addr;
  wire  mem_181_0_W0_clk;
  wire [7:0] mem_181_0_W0_data;
  wire  mem_181_0_W0_en;
  wire  mem_181_0_W0_mask;
  wire [25:0] mem_181_1_R0_addr;
  wire  mem_181_1_R0_clk;
  wire [7:0] mem_181_1_R0_data;
  wire  mem_181_1_R0_en;
  wire [25:0] mem_181_1_W0_addr;
  wire  mem_181_1_W0_clk;
  wire [7:0] mem_181_1_W0_data;
  wire  mem_181_1_W0_en;
  wire  mem_181_1_W0_mask;
  wire [25:0] mem_181_2_R0_addr;
  wire  mem_181_2_R0_clk;
  wire [7:0] mem_181_2_R0_data;
  wire  mem_181_2_R0_en;
  wire [25:0] mem_181_2_W0_addr;
  wire  mem_181_2_W0_clk;
  wire [7:0] mem_181_2_W0_data;
  wire  mem_181_2_W0_en;
  wire  mem_181_2_W0_mask;
  wire [25:0] mem_181_3_R0_addr;
  wire  mem_181_3_R0_clk;
  wire [7:0] mem_181_3_R0_data;
  wire  mem_181_3_R0_en;
  wire [25:0] mem_181_3_W0_addr;
  wire  mem_181_3_W0_clk;
  wire [7:0] mem_181_3_W0_data;
  wire  mem_181_3_W0_en;
  wire  mem_181_3_W0_mask;
  wire [25:0] mem_181_4_R0_addr;
  wire  mem_181_4_R0_clk;
  wire [7:0] mem_181_4_R0_data;
  wire  mem_181_4_R0_en;
  wire [25:0] mem_181_4_W0_addr;
  wire  mem_181_4_W0_clk;
  wire [7:0] mem_181_4_W0_data;
  wire  mem_181_4_W0_en;
  wire  mem_181_4_W0_mask;
  wire [25:0] mem_181_5_R0_addr;
  wire  mem_181_5_R0_clk;
  wire [7:0] mem_181_5_R0_data;
  wire  mem_181_5_R0_en;
  wire [25:0] mem_181_5_W0_addr;
  wire  mem_181_5_W0_clk;
  wire [7:0] mem_181_5_W0_data;
  wire  mem_181_5_W0_en;
  wire  mem_181_5_W0_mask;
  wire [25:0] mem_181_6_R0_addr;
  wire  mem_181_6_R0_clk;
  wire [7:0] mem_181_6_R0_data;
  wire  mem_181_6_R0_en;
  wire [25:0] mem_181_6_W0_addr;
  wire  mem_181_6_W0_clk;
  wire [7:0] mem_181_6_W0_data;
  wire  mem_181_6_W0_en;
  wire  mem_181_6_W0_mask;
  wire [25:0] mem_181_7_R0_addr;
  wire  mem_181_7_R0_clk;
  wire [7:0] mem_181_7_R0_data;
  wire  mem_181_7_R0_en;
  wire [25:0] mem_181_7_W0_addr;
  wire  mem_181_7_W0_clk;
  wire [7:0] mem_181_7_W0_data;
  wire  mem_181_7_W0_en;
  wire  mem_181_7_W0_mask;
  wire [25:0] mem_182_0_R0_addr;
  wire  mem_182_0_R0_clk;
  wire [7:0] mem_182_0_R0_data;
  wire  mem_182_0_R0_en;
  wire [25:0] mem_182_0_W0_addr;
  wire  mem_182_0_W0_clk;
  wire [7:0] mem_182_0_W0_data;
  wire  mem_182_0_W0_en;
  wire  mem_182_0_W0_mask;
  wire [25:0] mem_182_1_R0_addr;
  wire  mem_182_1_R0_clk;
  wire [7:0] mem_182_1_R0_data;
  wire  mem_182_1_R0_en;
  wire [25:0] mem_182_1_W0_addr;
  wire  mem_182_1_W0_clk;
  wire [7:0] mem_182_1_W0_data;
  wire  mem_182_1_W0_en;
  wire  mem_182_1_W0_mask;
  wire [25:0] mem_182_2_R0_addr;
  wire  mem_182_2_R0_clk;
  wire [7:0] mem_182_2_R0_data;
  wire  mem_182_2_R0_en;
  wire [25:0] mem_182_2_W0_addr;
  wire  mem_182_2_W0_clk;
  wire [7:0] mem_182_2_W0_data;
  wire  mem_182_2_W0_en;
  wire  mem_182_2_W0_mask;
  wire [25:0] mem_182_3_R0_addr;
  wire  mem_182_3_R0_clk;
  wire [7:0] mem_182_3_R0_data;
  wire  mem_182_3_R0_en;
  wire [25:0] mem_182_3_W0_addr;
  wire  mem_182_3_W0_clk;
  wire [7:0] mem_182_3_W0_data;
  wire  mem_182_3_W0_en;
  wire  mem_182_3_W0_mask;
  wire [25:0] mem_182_4_R0_addr;
  wire  mem_182_4_R0_clk;
  wire [7:0] mem_182_4_R0_data;
  wire  mem_182_4_R0_en;
  wire [25:0] mem_182_4_W0_addr;
  wire  mem_182_4_W0_clk;
  wire [7:0] mem_182_4_W0_data;
  wire  mem_182_4_W0_en;
  wire  mem_182_4_W0_mask;
  wire [25:0] mem_182_5_R0_addr;
  wire  mem_182_5_R0_clk;
  wire [7:0] mem_182_5_R0_data;
  wire  mem_182_5_R0_en;
  wire [25:0] mem_182_5_W0_addr;
  wire  mem_182_5_W0_clk;
  wire [7:0] mem_182_5_W0_data;
  wire  mem_182_5_W0_en;
  wire  mem_182_5_W0_mask;
  wire [25:0] mem_182_6_R0_addr;
  wire  mem_182_6_R0_clk;
  wire [7:0] mem_182_6_R0_data;
  wire  mem_182_6_R0_en;
  wire [25:0] mem_182_6_W0_addr;
  wire  mem_182_6_W0_clk;
  wire [7:0] mem_182_6_W0_data;
  wire  mem_182_6_W0_en;
  wire  mem_182_6_W0_mask;
  wire [25:0] mem_182_7_R0_addr;
  wire  mem_182_7_R0_clk;
  wire [7:0] mem_182_7_R0_data;
  wire  mem_182_7_R0_en;
  wire [25:0] mem_182_7_W0_addr;
  wire  mem_182_7_W0_clk;
  wire [7:0] mem_182_7_W0_data;
  wire  mem_182_7_W0_en;
  wire  mem_182_7_W0_mask;
  wire [25:0] mem_183_0_R0_addr;
  wire  mem_183_0_R0_clk;
  wire [7:0] mem_183_0_R0_data;
  wire  mem_183_0_R0_en;
  wire [25:0] mem_183_0_W0_addr;
  wire  mem_183_0_W0_clk;
  wire [7:0] mem_183_0_W0_data;
  wire  mem_183_0_W0_en;
  wire  mem_183_0_W0_mask;
  wire [25:0] mem_183_1_R0_addr;
  wire  mem_183_1_R0_clk;
  wire [7:0] mem_183_1_R0_data;
  wire  mem_183_1_R0_en;
  wire [25:0] mem_183_1_W0_addr;
  wire  mem_183_1_W0_clk;
  wire [7:0] mem_183_1_W0_data;
  wire  mem_183_1_W0_en;
  wire  mem_183_1_W0_mask;
  wire [25:0] mem_183_2_R0_addr;
  wire  mem_183_2_R0_clk;
  wire [7:0] mem_183_2_R0_data;
  wire  mem_183_2_R0_en;
  wire [25:0] mem_183_2_W0_addr;
  wire  mem_183_2_W0_clk;
  wire [7:0] mem_183_2_W0_data;
  wire  mem_183_2_W0_en;
  wire  mem_183_2_W0_mask;
  wire [25:0] mem_183_3_R0_addr;
  wire  mem_183_3_R0_clk;
  wire [7:0] mem_183_3_R0_data;
  wire  mem_183_3_R0_en;
  wire [25:0] mem_183_3_W0_addr;
  wire  mem_183_3_W0_clk;
  wire [7:0] mem_183_3_W0_data;
  wire  mem_183_3_W0_en;
  wire  mem_183_3_W0_mask;
  wire [25:0] mem_183_4_R0_addr;
  wire  mem_183_4_R0_clk;
  wire [7:0] mem_183_4_R0_data;
  wire  mem_183_4_R0_en;
  wire [25:0] mem_183_4_W0_addr;
  wire  mem_183_4_W0_clk;
  wire [7:0] mem_183_4_W0_data;
  wire  mem_183_4_W0_en;
  wire  mem_183_4_W0_mask;
  wire [25:0] mem_183_5_R0_addr;
  wire  mem_183_5_R0_clk;
  wire [7:0] mem_183_5_R0_data;
  wire  mem_183_5_R0_en;
  wire [25:0] mem_183_5_W0_addr;
  wire  mem_183_5_W0_clk;
  wire [7:0] mem_183_5_W0_data;
  wire  mem_183_5_W0_en;
  wire  mem_183_5_W0_mask;
  wire [25:0] mem_183_6_R0_addr;
  wire  mem_183_6_R0_clk;
  wire [7:0] mem_183_6_R0_data;
  wire  mem_183_6_R0_en;
  wire [25:0] mem_183_6_W0_addr;
  wire  mem_183_6_W0_clk;
  wire [7:0] mem_183_6_W0_data;
  wire  mem_183_6_W0_en;
  wire  mem_183_6_W0_mask;
  wire [25:0] mem_183_7_R0_addr;
  wire  mem_183_7_R0_clk;
  wire [7:0] mem_183_7_R0_data;
  wire  mem_183_7_R0_en;
  wire [25:0] mem_183_7_W0_addr;
  wire  mem_183_7_W0_clk;
  wire [7:0] mem_183_7_W0_data;
  wire  mem_183_7_W0_en;
  wire  mem_183_7_W0_mask;
  wire [25:0] mem_184_0_R0_addr;
  wire  mem_184_0_R0_clk;
  wire [7:0] mem_184_0_R0_data;
  wire  mem_184_0_R0_en;
  wire [25:0] mem_184_0_W0_addr;
  wire  mem_184_0_W0_clk;
  wire [7:0] mem_184_0_W0_data;
  wire  mem_184_0_W0_en;
  wire  mem_184_0_W0_mask;
  wire [25:0] mem_184_1_R0_addr;
  wire  mem_184_1_R0_clk;
  wire [7:0] mem_184_1_R0_data;
  wire  mem_184_1_R0_en;
  wire [25:0] mem_184_1_W0_addr;
  wire  mem_184_1_W0_clk;
  wire [7:0] mem_184_1_W0_data;
  wire  mem_184_1_W0_en;
  wire  mem_184_1_W0_mask;
  wire [25:0] mem_184_2_R0_addr;
  wire  mem_184_2_R0_clk;
  wire [7:0] mem_184_2_R0_data;
  wire  mem_184_2_R0_en;
  wire [25:0] mem_184_2_W0_addr;
  wire  mem_184_2_W0_clk;
  wire [7:0] mem_184_2_W0_data;
  wire  mem_184_2_W0_en;
  wire  mem_184_2_W0_mask;
  wire [25:0] mem_184_3_R0_addr;
  wire  mem_184_3_R0_clk;
  wire [7:0] mem_184_3_R0_data;
  wire  mem_184_3_R0_en;
  wire [25:0] mem_184_3_W0_addr;
  wire  mem_184_3_W0_clk;
  wire [7:0] mem_184_3_W0_data;
  wire  mem_184_3_W0_en;
  wire  mem_184_3_W0_mask;
  wire [25:0] mem_184_4_R0_addr;
  wire  mem_184_4_R0_clk;
  wire [7:0] mem_184_4_R0_data;
  wire  mem_184_4_R0_en;
  wire [25:0] mem_184_4_W0_addr;
  wire  mem_184_4_W0_clk;
  wire [7:0] mem_184_4_W0_data;
  wire  mem_184_4_W0_en;
  wire  mem_184_4_W0_mask;
  wire [25:0] mem_184_5_R0_addr;
  wire  mem_184_5_R0_clk;
  wire [7:0] mem_184_5_R0_data;
  wire  mem_184_5_R0_en;
  wire [25:0] mem_184_5_W0_addr;
  wire  mem_184_5_W0_clk;
  wire [7:0] mem_184_5_W0_data;
  wire  mem_184_5_W0_en;
  wire  mem_184_5_W0_mask;
  wire [25:0] mem_184_6_R0_addr;
  wire  mem_184_6_R0_clk;
  wire [7:0] mem_184_6_R0_data;
  wire  mem_184_6_R0_en;
  wire [25:0] mem_184_6_W0_addr;
  wire  mem_184_6_W0_clk;
  wire [7:0] mem_184_6_W0_data;
  wire  mem_184_6_W0_en;
  wire  mem_184_6_W0_mask;
  wire [25:0] mem_184_7_R0_addr;
  wire  mem_184_7_R0_clk;
  wire [7:0] mem_184_7_R0_data;
  wire  mem_184_7_R0_en;
  wire [25:0] mem_184_7_W0_addr;
  wire  mem_184_7_W0_clk;
  wire [7:0] mem_184_7_W0_data;
  wire  mem_184_7_W0_en;
  wire  mem_184_7_W0_mask;
  wire [25:0] mem_185_0_R0_addr;
  wire  mem_185_0_R0_clk;
  wire [7:0] mem_185_0_R0_data;
  wire  mem_185_0_R0_en;
  wire [25:0] mem_185_0_W0_addr;
  wire  mem_185_0_W0_clk;
  wire [7:0] mem_185_0_W0_data;
  wire  mem_185_0_W0_en;
  wire  mem_185_0_W0_mask;
  wire [25:0] mem_185_1_R0_addr;
  wire  mem_185_1_R0_clk;
  wire [7:0] mem_185_1_R0_data;
  wire  mem_185_1_R0_en;
  wire [25:0] mem_185_1_W0_addr;
  wire  mem_185_1_W0_clk;
  wire [7:0] mem_185_1_W0_data;
  wire  mem_185_1_W0_en;
  wire  mem_185_1_W0_mask;
  wire [25:0] mem_185_2_R0_addr;
  wire  mem_185_2_R0_clk;
  wire [7:0] mem_185_2_R0_data;
  wire  mem_185_2_R0_en;
  wire [25:0] mem_185_2_W0_addr;
  wire  mem_185_2_W0_clk;
  wire [7:0] mem_185_2_W0_data;
  wire  mem_185_2_W0_en;
  wire  mem_185_2_W0_mask;
  wire [25:0] mem_185_3_R0_addr;
  wire  mem_185_3_R0_clk;
  wire [7:0] mem_185_3_R0_data;
  wire  mem_185_3_R0_en;
  wire [25:0] mem_185_3_W0_addr;
  wire  mem_185_3_W0_clk;
  wire [7:0] mem_185_3_W0_data;
  wire  mem_185_3_W0_en;
  wire  mem_185_3_W0_mask;
  wire [25:0] mem_185_4_R0_addr;
  wire  mem_185_4_R0_clk;
  wire [7:0] mem_185_4_R0_data;
  wire  mem_185_4_R0_en;
  wire [25:0] mem_185_4_W0_addr;
  wire  mem_185_4_W0_clk;
  wire [7:0] mem_185_4_W0_data;
  wire  mem_185_4_W0_en;
  wire  mem_185_4_W0_mask;
  wire [25:0] mem_185_5_R0_addr;
  wire  mem_185_5_R0_clk;
  wire [7:0] mem_185_5_R0_data;
  wire  mem_185_5_R0_en;
  wire [25:0] mem_185_5_W0_addr;
  wire  mem_185_5_W0_clk;
  wire [7:0] mem_185_5_W0_data;
  wire  mem_185_5_W0_en;
  wire  mem_185_5_W0_mask;
  wire [25:0] mem_185_6_R0_addr;
  wire  mem_185_6_R0_clk;
  wire [7:0] mem_185_6_R0_data;
  wire  mem_185_6_R0_en;
  wire [25:0] mem_185_6_W0_addr;
  wire  mem_185_6_W0_clk;
  wire [7:0] mem_185_6_W0_data;
  wire  mem_185_6_W0_en;
  wire  mem_185_6_W0_mask;
  wire [25:0] mem_185_7_R0_addr;
  wire  mem_185_7_R0_clk;
  wire [7:0] mem_185_7_R0_data;
  wire  mem_185_7_R0_en;
  wire [25:0] mem_185_7_W0_addr;
  wire  mem_185_7_W0_clk;
  wire [7:0] mem_185_7_W0_data;
  wire  mem_185_7_W0_en;
  wire  mem_185_7_W0_mask;
  wire [25:0] mem_186_0_R0_addr;
  wire  mem_186_0_R0_clk;
  wire [7:0] mem_186_0_R0_data;
  wire  mem_186_0_R0_en;
  wire [25:0] mem_186_0_W0_addr;
  wire  mem_186_0_W0_clk;
  wire [7:0] mem_186_0_W0_data;
  wire  mem_186_0_W0_en;
  wire  mem_186_0_W0_mask;
  wire [25:0] mem_186_1_R0_addr;
  wire  mem_186_1_R0_clk;
  wire [7:0] mem_186_1_R0_data;
  wire  mem_186_1_R0_en;
  wire [25:0] mem_186_1_W0_addr;
  wire  mem_186_1_W0_clk;
  wire [7:0] mem_186_1_W0_data;
  wire  mem_186_1_W0_en;
  wire  mem_186_1_W0_mask;
  wire [25:0] mem_186_2_R0_addr;
  wire  mem_186_2_R0_clk;
  wire [7:0] mem_186_2_R0_data;
  wire  mem_186_2_R0_en;
  wire [25:0] mem_186_2_W0_addr;
  wire  mem_186_2_W0_clk;
  wire [7:0] mem_186_2_W0_data;
  wire  mem_186_2_W0_en;
  wire  mem_186_2_W0_mask;
  wire [25:0] mem_186_3_R0_addr;
  wire  mem_186_3_R0_clk;
  wire [7:0] mem_186_3_R0_data;
  wire  mem_186_3_R0_en;
  wire [25:0] mem_186_3_W0_addr;
  wire  mem_186_3_W0_clk;
  wire [7:0] mem_186_3_W0_data;
  wire  mem_186_3_W0_en;
  wire  mem_186_3_W0_mask;
  wire [25:0] mem_186_4_R0_addr;
  wire  mem_186_4_R0_clk;
  wire [7:0] mem_186_4_R0_data;
  wire  mem_186_4_R0_en;
  wire [25:0] mem_186_4_W0_addr;
  wire  mem_186_4_W0_clk;
  wire [7:0] mem_186_4_W0_data;
  wire  mem_186_4_W0_en;
  wire  mem_186_4_W0_mask;
  wire [25:0] mem_186_5_R0_addr;
  wire  mem_186_5_R0_clk;
  wire [7:0] mem_186_5_R0_data;
  wire  mem_186_5_R0_en;
  wire [25:0] mem_186_5_W0_addr;
  wire  mem_186_5_W0_clk;
  wire [7:0] mem_186_5_W0_data;
  wire  mem_186_5_W0_en;
  wire  mem_186_5_W0_mask;
  wire [25:0] mem_186_6_R0_addr;
  wire  mem_186_6_R0_clk;
  wire [7:0] mem_186_6_R0_data;
  wire  mem_186_6_R0_en;
  wire [25:0] mem_186_6_W0_addr;
  wire  mem_186_6_W0_clk;
  wire [7:0] mem_186_6_W0_data;
  wire  mem_186_6_W0_en;
  wire  mem_186_6_W0_mask;
  wire [25:0] mem_186_7_R0_addr;
  wire  mem_186_7_R0_clk;
  wire [7:0] mem_186_7_R0_data;
  wire  mem_186_7_R0_en;
  wire [25:0] mem_186_7_W0_addr;
  wire  mem_186_7_W0_clk;
  wire [7:0] mem_186_7_W0_data;
  wire  mem_186_7_W0_en;
  wire  mem_186_7_W0_mask;
  wire [25:0] mem_187_0_R0_addr;
  wire  mem_187_0_R0_clk;
  wire [7:0] mem_187_0_R0_data;
  wire  mem_187_0_R0_en;
  wire [25:0] mem_187_0_W0_addr;
  wire  mem_187_0_W0_clk;
  wire [7:0] mem_187_0_W0_data;
  wire  mem_187_0_W0_en;
  wire  mem_187_0_W0_mask;
  wire [25:0] mem_187_1_R0_addr;
  wire  mem_187_1_R0_clk;
  wire [7:0] mem_187_1_R0_data;
  wire  mem_187_1_R0_en;
  wire [25:0] mem_187_1_W0_addr;
  wire  mem_187_1_W0_clk;
  wire [7:0] mem_187_1_W0_data;
  wire  mem_187_1_W0_en;
  wire  mem_187_1_W0_mask;
  wire [25:0] mem_187_2_R0_addr;
  wire  mem_187_2_R0_clk;
  wire [7:0] mem_187_2_R0_data;
  wire  mem_187_2_R0_en;
  wire [25:0] mem_187_2_W0_addr;
  wire  mem_187_2_W0_clk;
  wire [7:0] mem_187_2_W0_data;
  wire  mem_187_2_W0_en;
  wire  mem_187_2_W0_mask;
  wire [25:0] mem_187_3_R0_addr;
  wire  mem_187_3_R0_clk;
  wire [7:0] mem_187_3_R0_data;
  wire  mem_187_3_R0_en;
  wire [25:0] mem_187_3_W0_addr;
  wire  mem_187_3_W0_clk;
  wire [7:0] mem_187_3_W0_data;
  wire  mem_187_3_W0_en;
  wire  mem_187_3_W0_mask;
  wire [25:0] mem_187_4_R0_addr;
  wire  mem_187_4_R0_clk;
  wire [7:0] mem_187_4_R0_data;
  wire  mem_187_4_R0_en;
  wire [25:0] mem_187_4_W0_addr;
  wire  mem_187_4_W0_clk;
  wire [7:0] mem_187_4_W0_data;
  wire  mem_187_4_W0_en;
  wire  mem_187_4_W0_mask;
  wire [25:0] mem_187_5_R0_addr;
  wire  mem_187_5_R0_clk;
  wire [7:0] mem_187_5_R0_data;
  wire  mem_187_5_R0_en;
  wire [25:0] mem_187_5_W0_addr;
  wire  mem_187_5_W0_clk;
  wire [7:0] mem_187_5_W0_data;
  wire  mem_187_5_W0_en;
  wire  mem_187_5_W0_mask;
  wire [25:0] mem_187_6_R0_addr;
  wire  mem_187_6_R0_clk;
  wire [7:0] mem_187_6_R0_data;
  wire  mem_187_6_R0_en;
  wire [25:0] mem_187_6_W0_addr;
  wire  mem_187_6_W0_clk;
  wire [7:0] mem_187_6_W0_data;
  wire  mem_187_6_W0_en;
  wire  mem_187_6_W0_mask;
  wire [25:0] mem_187_7_R0_addr;
  wire  mem_187_7_R0_clk;
  wire [7:0] mem_187_7_R0_data;
  wire  mem_187_7_R0_en;
  wire [25:0] mem_187_7_W0_addr;
  wire  mem_187_7_W0_clk;
  wire [7:0] mem_187_7_W0_data;
  wire  mem_187_7_W0_en;
  wire  mem_187_7_W0_mask;
  wire [25:0] mem_188_0_R0_addr;
  wire  mem_188_0_R0_clk;
  wire [7:0] mem_188_0_R0_data;
  wire  mem_188_0_R0_en;
  wire [25:0] mem_188_0_W0_addr;
  wire  mem_188_0_W0_clk;
  wire [7:0] mem_188_0_W0_data;
  wire  mem_188_0_W0_en;
  wire  mem_188_0_W0_mask;
  wire [25:0] mem_188_1_R0_addr;
  wire  mem_188_1_R0_clk;
  wire [7:0] mem_188_1_R0_data;
  wire  mem_188_1_R0_en;
  wire [25:0] mem_188_1_W0_addr;
  wire  mem_188_1_W0_clk;
  wire [7:0] mem_188_1_W0_data;
  wire  mem_188_1_W0_en;
  wire  mem_188_1_W0_mask;
  wire [25:0] mem_188_2_R0_addr;
  wire  mem_188_2_R0_clk;
  wire [7:0] mem_188_2_R0_data;
  wire  mem_188_2_R0_en;
  wire [25:0] mem_188_2_W0_addr;
  wire  mem_188_2_W0_clk;
  wire [7:0] mem_188_2_W0_data;
  wire  mem_188_2_W0_en;
  wire  mem_188_2_W0_mask;
  wire [25:0] mem_188_3_R0_addr;
  wire  mem_188_3_R0_clk;
  wire [7:0] mem_188_3_R0_data;
  wire  mem_188_3_R0_en;
  wire [25:0] mem_188_3_W0_addr;
  wire  mem_188_3_W0_clk;
  wire [7:0] mem_188_3_W0_data;
  wire  mem_188_3_W0_en;
  wire  mem_188_3_W0_mask;
  wire [25:0] mem_188_4_R0_addr;
  wire  mem_188_4_R0_clk;
  wire [7:0] mem_188_4_R0_data;
  wire  mem_188_4_R0_en;
  wire [25:0] mem_188_4_W0_addr;
  wire  mem_188_4_W0_clk;
  wire [7:0] mem_188_4_W0_data;
  wire  mem_188_4_W0_en;
  wire  mem_188_4_W0_mask;
  wire [25:0] mem_188_5_R0_addr;
  wire  mem_188_5_R0_clk;
  wire [7:0] mem_188_5_R0_data;
  wire  mem_188_5_R0_en;
  wire [25:0] mem_188_5_W0_addr;
  wire  mem_188_5_W0_clk;
  wire [7:0] mem_188_5_W0_data;
  wire  mem_188_5_W0_en;
  wire  mem_188_5_W0_mask;
  wire [25:0] mem_188_6_R0_addr;
  wire  mem_188_6_R0_clk;
  wire [7:0] mem_188_6_R0_data;
  wire  mem_188_6_R0_en;
  wire [25:0] mem_188_6_W0_addr;
  wire  mem_188_6_W0_clk;
  wire [7:0] mem_188_6_W0_data;
  wire  mem_188_6_W0_en;
  wire  mem_188_6_W0_mask;
  wire [25:0] mem_188_7_R0_addr;
  wire  mem_188_7_R0_clk;
  wire [7:0] mem_188_7_R0_data;
  wire  mem_188_7_R0_en;
  wire [25:0] mem_188_7_W0_addr;
  wire  mem_188_7_W0_clk;
  wire [7:0] mem_188_7_W0_data;
  wire  mem_188_7_W0_en;
  wire  mem_188_7_W0_mask;
  wire [25:0] mem_189_0_R0_addr;
  wire  mem_189_0_R0_clk;
  wire [7:0] mem_189_0_R0_data;
  wire  mem_189_0_R0_en;
  wire [25:0] mem_189_0_W0_addr;
  wire  mem_189_0_W0_clk;
  wire [7:0] mem_189_0_W0_data;
  wire  mem_189_0_W0_en;
  wire  mem_189_0_W0_mask;
  wire [25:0] mem_189_1_R0_addr;
  wire  mem_189_1_R0_clk;
  wire [7:0] mem_189_1_R0_data;
  wire  mem_189_1_R0_en;
  wire [25:0] mem_189_1_W0_addr;
  wire  mem_189_1_W0_clk;
  wire [7:0] mem_189_1_W0_data;
  wire  mem_189_1_W0_en;
  wire  mem_189_1_W0_mask;
  wire [25:0] mem_189_2_R0_addr;
  wire  mem_189_2_R0_clk;
  wire [7:0] mem_189_2_R0_data;
  wire  mem_189_2_R0_en;
  wire [25:0] mem_189_2_W0_addr;
  wire  mem_189_2_W0_clk;
  wire [7:0] mem_189_2_W0_data;
  wire  mem_189_2_W0_en;
  wire  mem_189_2_W0_mask;
  wire [25:0] mem_189_3_R0_addr;
  wire  mem_189_3_R0_clk;
  wire [7:0] mem_189_3_R0_data;
  wire  mem_189_3_R0_en;
  wire [25:0] mem_189_3_W0_addr;
  wire  mem_189_3_W0_clk;
  wire [7:0] mem_189_3_W0_data;
  wire  mem_189_3_W0_en;
  wire  mem_189_3_W0_mask;
  wire [25:0] mem_189_4_R0_addr;
  wire  mem_189_4_R0_clk;
  wire [7:0] mem_189_4_R0_data;
  wire  mem_189_4_R0_en;
  wire [25:0] mem_189_4_W0_addr;
  wire  mem_189_4_W0_clk;
  wire [7:0] mem_189_4_W0_data;
  wire  mem_189_4_W0_en;
  wire  mem_189_4_W0_mask;
  wire [25:0] mem_189_5_R0_addr;
  wire  mem_189_5_R0_clk;
  wire [7:0] mem_189_5_R0_data;
  wire  mem_189_5_R0_en;
  wire [25:0] mem_189_5_W0_addr;
  wire  mem_189_5_W0_clk;
  wire [7:0] mem_189_5_W0_data;
  wire  mem_189_5_W0_en;
  wire  mem_189_5_W0_mask;
  wire [25:0] mem_189_6_R0_addr;
  wire  mem_189_6_R0_clk;
  wire [7:0] mem_189_6_R0_data;
  wire  mem_189_6_R0_en;
  wire [25:0] mem_189_6_W0_addr;
  wire  mem_189_6_W0_clk;
  wire [7:0] mem_189_6_W0_data;
  wire  mem_189_6_W0_en;
  wire  mem_189_6_W0_mask;
  wire [25:0] mem_189_7_R0_addr;
  wire  mem_189_7_R0_clk;
  wire [7:0] mem_189_7_R0_data;
  wire  mem_189_7_R0_en;
  wire [25:0] mem_189_7_W0_addr;
  wire  mem_189_7_W0_clk;
  wire [7:0] mem_189_7_W0_data;
  wire  mem_189_7_W0_en;
  wire  mem_189_7_W0_mask;
  wire [25:0] mem_190_0_R0_addr;
  wire  mem_190_0_R0_clk;
  wire [7:0] mem_190_0_R0_data;
  wire  mem_190_0_R0_en;
  wire [25:0] mem_190_0_W0_addr;
  wire  mem_190_0_W0_clk;
  wire [7:0] mem_190_0_W0_data;
  wire  mem_190_0_W0_en;
  wire  mem_190_0_W0_mask;
  wire [25:0] mem_190_1_R0_addr;
  wire  mem_190_1_R0_clk;
  wire [7:0] mem_190_1_R0_data;
  wire  mem_190_1_R0_en;
  wire [25:0] mem_190_1_W0_addr;
  wire  mem_190_1_W0_clk;
  wire [7:0] mem_190_1_W0_data;
  wire  mem_190_1_W0_en;
  wire  mem_190_1_W0_mask;
  wire [25:0] mem_190_2_R0_addr;
  wire  mem_190_2_R0_clk;
  wire [7:0] mem_190_2_R0_data;
  wire  mem_190_2_R0_en;
  wire [25:0] mem_190_2_W0_addr;
  wire  mem_190_2_W0_clk;
  wire [7:0] mem_190_2_W0_data;
  wire  mem_190_2_W0_en;
  wire  mem_190_2_W0_mask;
  wire [25:0] mem_190_3_R0_addr;
  wire  mem_190_3_R0_clk;
  wire [7:0] mem_190_3_R0_data;
  wire  mem_190_3_R0_en;
  wire [25:0] mem_190_3_W0_addr;
  wire  mem_190_3_W0_clk;
  wire [7:0] mem_190_3_W0_data;
  wire  mem_190_3_W0_en;
  wire  mem_190_3_W0_mask;
  wire [25:0] mem_190_4_R0_addr;
  wire  mem_190_4_R0_clk;
  wire [7:0] mem_190_4_R0_data;
  wire  mem_190_4_R0_en;
  wire [25:0] mem_190_4_W0_addr;
  wire  mem_190_4_W0_clk;
  wire [7:0] mem_190_4_W0_data;
  wire  mem_190_4_W0_en;
  wire  mem_190_4_W0_mask;
  wire [25:0] mem_190_5_R0_addr;
  wire  mem_190_5_R0_clk;
  wire [7:0] mem_190_5_R0_data;
  wire  mem_190_5_R0_en;
  wire [25:0] mem_190_5_W0_addr;
  wire  mem_190_5_W0_clk;
  wire [7:0] mem_190_5_W0_data;
  wire  mem_190_5_W0_en;
  wire  mem_190_5_W0_mask;
  wire [25:0] mem_190_6_R0_addr;
  wire  mem_190_6_R0_clk;
  wire [7:0] mem_190_6_R0_data;
  wire  mem_190_6_R0_en;
  wire [25:0] mem_190_6_W0_addr;
  wire  mem_190_6_W0_clk;
  wire [7:0] mem_190_6_W0_data;
  wire  mem_190_6_W0_en;
  wire  mem_190_6_W0_mask;
  wire [25:0] mem_190_7_R0_addr;
  wire  mem_190_7_R0_clk;
  wire [7:0] mem_190_7_R0_data;
  wire  mem_190_7_R0_en;
  wire [25:0] mem_190_7_W0_addr;
  wire  mem_190_7_W0_clk;
  wire [7:0] mem_190_7_W0_data;
  wire  mem_190_7_W0_en;
  wire  mem_190_7_W0_mask;
  wire [25:0] mem_191_0_R0_addr;
  wire  mem_191_0_R0_clk;
  wire [7:0] mem_191_0_R0_data;
  wire  mem_191_0_R0_en;
  wire [25:0] mem_191_0_W0_addr;
  wire  mem_191_0_W0_clk;
  wire [7:0] mem_191_0_W0_data;
  wire  mem_191_0_W0_en;
  wire  mem_191_0_W0_mask;
  wire [25:0] mem_191_1_R0_addr;
  wire  mem_191_1_R0_clk;
  wire [7:0] mem_191_1_R0_data;
  wire  mem_191_1_R0_en;
  wire [25:0] mem_191_1_W0_addr;
  wire  mem_191_1_W0_clk;
  wire [7:0] mem_191_1_W0_data;
  wire  mem_191_1_W0_en;
  wire  mem_191_1_W0_mask;
  wire [25:0] mem_191_2_R0_addr;
  wire  mem_191_2_R0_clk;
  wire [7:0] mem_191_2_R0_data;
  wire  mem_191_2_R0_en;
  wire [25:0] mem_191_2_W0_addr;
  wire  mem_191_2_W0_clk;
  wire [7:0] mem_191_2_W0_data;
  wire  mem_191_2_W0_en;
  wire  mem_191_2_W0_mask;
  wire [25:0] mem_191_3_R0_addr;
  wire  mem_191_3_R0_clk;
  wire [7:0] mem_191_3_R0_data;
  wire  mem_191_3_R0_en;
  wire [25:0] mem_191_3_W0_addr;
  wire  mem_191_3_W0_clk;
  wire [7:0] mem_191_3_W0_data;
  wire  mem_191_3_W0_en;
  wire  mem_191_3_W0_mask;
  wire [25:0] mem_191_4_R0_addr;
  wire  mem_191_4_R0_clk;
  wire [7:0] mem_191_4_R0_data;
  wire  mem_191_4_R0_en;
  wire [25:0] mem_191_4_W0_addr;
  wire  mem_191_4_W0_clk;
  wire [7:0] mem_191_4_W0_data;
  wire  mem_191_4_W0_en;
  wire  mem_191_4_W0_mask;
  wire [25:0] mem_191_5_R0_addr;
  wire  mem_191_5_R0_clk;
  wire [7:0] mem_191_5_R0_data;
  wire  mem_191_5_R0_en;
  wire [25:0] mem_191_5_W0_addr;
  wire  mem_191_5_W0_clk;
  wire [7:0] mem_191_5_W0_data;
  wire  mem_191_5_W0_en;
  wire  mem_191_5_W0_mask;
  wire [25:0] mem_191_6_R0_addr;
  wire  mem_191_6_R0_clk;
  wire [7:0] mem_191_6_R0_data;
  wire  mem_191_6_R0_en;
  wire [25:0] mem_191_6_W0_addr;
  wire  mem_191_6_W0_clk;
  wire [7:0] mem_191_6_W0_data;
  wire  mem_191_6_W0_en;
  wire  mem_191_6_W0_mask;
  wire [25:0] mem_191_7_R0_addr;
  wire  mem_191_7_R0_clk;
  wire [7:0] mem_191_7_R0_data;
  wire  mem_191_7_R0_en;
  wire [25:0] mem_191_7_W0_addr;
  wire  mem_191_7_W0_clk;
  wire [7:0] mem_191_7_W0_data;
  wire  mem_191_7_W0_en;
  wire  mem_191_7_W0_mask;
  wire [25:0] mem_192_0_R0_addr;
  wire  mem_192_0_R0_clk;
  wire [7:0] mem_192_0_R0_data;
  wire  mem_192_0_R0_en;
  wire [25:0] mem_192_0_W0_addr;
  wire  mem_192_0_W0_clk;
  wire [7:0] mem_192_0_W0_data;
  wire  mem_192_0_W0_en;
  wire  mem_192_0_W0_mask;
  wire [25:0] mem_192_1_R0_addr;
  wire  mem_192_1_R0_clk;
  wire [7:0] mem_192_1_R0_data;
  wire  mem_192_1_R0_en;
  wire [25:0] mem_192_1_W0_addr;
  wire  mem_192_1_W0_clk;
  wire [7:0] mem_192_1_W0_data;
  wire  mem_192_1_W0_en;
  wire  mem_192_1_W0_mask;
  wire [25:0] mem_192_2_R0_addr;
  wire  mem_192_2_R0_clk;
  wire [7:0] mem_192_2_R0_data;
  wire  mem_192_2_R0_en;
  wire [25:0] mem_192_2_W0_addr;
  wire  mem_192_2_W0_clk;
  wire [7:0] mem_192_2_W0_data;
  wire  mem_192_2_W0_en;
  wire  mem_192_2_W0_mask;
  wire [25:0] mem_192_3_R0_addr;
  wire  mem_192_3_R0_clk;
  wire [7:0] mem_192_3_R0_data;
  wire  mem_192_3_R0_en;
  wire [25:0] mem_192_3_W0_addr;
  wire  mem_192_3_W0_clk;
  wire [7:0] mem_192_3_W0_data;
  wire  mem_192_3_W0_en;
  wire  mem_192_3_W0_mask;
  wire [25:0] mem_192_4_R0_addr;
  wire  mem_192_4_R0_clk;
  wire [7:0] mem_192_4_R0_data;
  wire  mem_192_4_R0_en;
  wire [25:0] mem_192_4_W0_addr;
  wire  mem_192_4_W0_clk;
  wire [7:0] mem_192_4_W0_data;
  wire  mem_192_4_W0_en;
  wire  mem_192_4_W0_mask;
  wire [25:0] mem_192_5_R0_addr;
  wire  mem_192_5_R0_clk;
  wire [7:0] mem_192_5_R0_data;
  wire  mem_192_5_R0_en;
  wire [25:0] mem_192_5_W0_addr;
  wire  mem_192_5_W0_clk;
  wire [7:0] mem_192_5_W0_data;
  wire  mem_192_5_W0_en;
  wire  mem_192_5_W0_mask;
  wire [25:0] mem_192_6_R0_addr;
  wire  mem_192_6_R0_clk;
  wire [7:0] mem_192_6_R0_data;
  wire  mem_192_6_R0_en;
  wire [25:0] mem_192_6_W0_addr;
  wire  mem_192_6_W0_clk;
  wire [7:0] mem_192_6_W0_data;
  wire  mem_192_6_W0_en;
  wire  mem_192_6_W0_mask;
  wire [25:0] mem_192_7_R0_addr;
  wire  mem_192_7_R0_clk;
  wire [7:0] mem_192_7_R0_data;
  wire  mem_192_7_R0_en;
  wire [25:0] mem_192_7_W0_addr;
  wire  mem_192_7_W0_clk;
  wire [7:0] mem_192_7_W0_data;
  wire  mem_192_7_W0_en;
  wire  mem_192_7_W0_mask;
  wire [25:0] mem_193_0_R0_addr;
  wire  mem_193_0_R0_clk;
  wire [7:0] mem_193_0_R0_data;
  wire  mem_193_0_R0_en;
  wire [25:0] mem_193_0_W0_addr;
  wire  mem_193_0_W0_clk;
  wire [7:0] mem_193_0_W0_data;
  wire  mem_193_0_W0_en;
  wire  mem_193_0_W0_mask;
  wire [25:0] mem_193_1_R0_addr;
  wire  mem_193_1_R0_clk;
  wire [7:0] mem_193_1_R0_data;
  wire  mem_193_1_R0_en;
  wire [25:0] mem_193_1_W0_addr;
  wire  mem_193_1_W0_clk;
  wire [7:0] mem_193_1_W0_data;
  wire  mem_193_1_W0_en;
  wire  mem_193_1_W0_mask;
  wire [25:0] mem_193_2_R0_addr;
  wire  mem_193_2_R0_clk;
  wire [7:0] mem_193_2_R0_data;
  wire  mem_193_2_R0_en;
  wire [25:0] mem_193_2_W0_addr;
  wire  mem_193_2_W0_clk;
  wire [7:0] mem_193_2_W0_data;
  wire  mem_193_2_W0_en;
  wire  mem_193_2_W0_mask;
  wire [25:0] mem_193_3_R0_addr;
  wire  mem_193_3_R0_clk;
  wire [7:0] mem_193_3_R0_data;
  wire  mem_193_3_R0_en;
  wire [25:0] mem_193_3_W0_addr;
  wire  mem_193_3_W0_clk;
  wire [7:0] mem_193_3_W0_data;
  wire  mem_193_3_W0_en;
  wire  mem_193_3_W0_mask;
  wire [25:0] mem_193_4_R0_addr;
  wire  mem_193_4_R0_clk;
  wire [7:0] mem_193_4_R0_data;
  wire  mem_193_4_R0_en;
  wire [25:0] mem_193_4_W0_addr;
  wire  mem_193_4_W0_clk;
  wire [7:0] mem_193_4_W0_data;
  wire  mem_193_4_W0_en;
  wire  mem_193_4_W0_mask;
  wire [25:0] mem_193_5_R0_addr;
  wire  mem_193_5_R0_clk;
  wire [7:0] mem_193_5_R0_data;
  wire  mem_193_5_R0_en;
  wire [25:0] mem_193_5_W0_addr;
  wire  mem_193_5_W0_clk;
  wire [7:0] mem_193_5_W0_data;
  wire  mem_193_5_W0_en;
  wire  mem_193_5_W0_mask;
  wire [25:0] mem_193_6_R0_addr;
  wire  mem_193_6_R0_clk;
  wire [7:0] mem_193_6_R0_data;
  wire  mem_193_6_R0_en;
  wire [25:0] mem_193_6_W0_addr;
  wire  mem_193_6_W0_clk;
  wire [7:0] mem_193_6_W0_data;
  wire  mem_193_6_W0_en;
  wire  mem_193_6_W0_mask;
  wire [25:0] mem_193_7_R0_addr;
  wire  mem_193_7_R0_clk;
  wire [7:0] mem_193_7_R0_data;
  wire  mem_193_7_R0_en;
  wire [25:0] mem_193_7_W0_addr;
  wire  mem_193_7_W0_clk;
  wire [7:0] mem_193_7_W0_data;
  wire  mem_193_7_W0_en;
  wire  mem_193_7_W0_mask;
  wire [25:0] mem_194_0_R0_addr;
  wire  mem_194_0_R0_clk;
  wire [7:0] mem_194_0_R0_data;
  wire  mem_194_0_R0_en;
  wire [25:0] mem_194_0_W0_addr;
  wire  mem_194_0_W0_clk;
  wire [7:0] mem_194_0_W0_data;
  wire  mem_194_0_W0_en;
  wire  mem_194_0_W0_mask;
  wire [25:0] mem_194_1_R0_addr;
  wire  mem_194_1_R0_clk;
  wire [7:0] mem_194_1_R0_data;
  wire  mem_194_1_R0_en;
  wire [25:0] mem_194_1_W0_addr;
  wire  mem_194_1_W0_clk;
  wire [7:0] mem_194_1_W0_data;
  wire  mem_194_1_W0_en;
  wire  mem_194_1_W0_mask;
  wire [25:0] mem_194_2_R0_addr;
  wire  mem_194_2_R0_clk;
  wire [7:0] mem_194_2_R0_data;
  wire  mem_194_2_R0_en;
  wire [25:0] mem_194_2_W0_addr;
  wire  mem_194_2_W0_clk;
  wire [7:0] mem_194_2_W0_data;
  wire  mem_194_2_W0_en;
  wire  mem_194_2_W0_mask;
  wire [25:0] mem_194_3_R0_addr;
  wire  mem_194_3_R0_clk;
  wire [7:0] mem_194_3_R0_data;
  wire  mem_194_3_R0_en;
  wire [25:0] mem_194_3_W0_addr;
  wire  mem_194_3_W0_clk;
  wire [7:0] mem_194_3_W0_data;
  wire  mem_194_3_W0_en;
  wire  mem_194_3_W0_mask;
  wire [25:0] mem_194_4_R0_addr;
  wire  mem_194_4_R0_clk;
  wire [7:0] mem_194_4_R0_data;
  wire  mem_194_4_R0_en;
  wire [25:0] mem_194_4_W0_addr;
  wire  mem_194_4_W0_clk;
  wire [7:0] mem_194_4_W0_data;
  wire  mem_194_4_W0_en;
  wire  mem_194_4_W0_mask;
  wire [25:0] mem_194_5_R0_addr;
  wire  mem_194_5_R0_clk;
  wire [7:0] mem_194_5_R0_data;
  wire  mem_194_5_R0_en;
  wire [25:0] mem_194_5_W0_addr;
  wire  mem_194_5_W0_clk;
  wire [7:0] mem_194_5_W0_data;
  wire  mem_194_5_W0_en;
  wire  mem_194_5_W0_mask;
  wire [25:0] mem_194_6_R0_addr;
  wire  mem_194_6_R0_clk;
  wire [7:0] mem_194_6_R0_data;
  wire  mem_194_6_R0_en;
  wire [25:0] mem_194_6_W0_addr;
  wire  mem_194_6_W0_clk;
  wire [7:0] mem_194_6_W0_data;
  wire  mem_194_6_W0_en;
  wire  mem_194_6_W0_mask;
  wire [25:0] mem_194_7_R0_addr;
  wire  mem_194_7_R0_clk;
  wire [7:0] mem_194_7_R0_data;
  wire  mem_194_7_R0_en;
  wire [25:0] mem_194_7_W0_addr;
  wire  mem_194_7_W0_clk;
  wire [7:0] mem_194_7_W0_data;
  wire  mem_194_7_W0_en;
  wire  mem_194_7_W0_mask;
  wire [25:0] mem_195_0_R0_addr;
  wire  mem_195_0_R0_clk;
  wire [7:0] mem_195_0_R0_data;
  wire  mem_195_0_R0_en;
  wire [25:0] mem_195_0_W0_addr;
  wire  mem_195_0_W0_clk;
  wire [7:0] mem_195_0_W0_data;
  wire  mem_195_0_W0_en;
  wire  mem_195_0_W0_mask;
  wire [25:0] mem_195_1_R0_addr;
  wire  mem_195_1_R0_clk;
  wire [7:0] mem_195_1_R0_data;
  wire  mem_195_1_R0_en;
  wire [25:0] mem_195_1_W0_addr;
  wire  mem_195_1_W0_clk;
  wire [7:0] mem_195_1_W0_data;
  wire  mem_195_1_W0_en;
  wire  mem_195_1_W0_mask;
  wire [25:0] mem_195_2_R0_addr;
  wire  mem_195_2_R0_clk;
  wire [7:0] mem_195_2_R0_data;
  wire  mem_195_2_R0_en;
  wire [25:0] mem_195_2_W0_addr;
  wire  mem_195_2_W0_clk;
  wire [7:0] mem_195_2_W0_data;
  wire  mem_195_2_W0_en;
  wire  mem_195_2_W0_mask;
  wire [25:0] mem_195_3_R0_addr;
  wire  mem_195_3_R0_clk;
  wire [7:0] mem_195_3_R0_data;
  wire  mem_195_3_R0_en;
  wire [25:0] mem_195_3_W0_addr;
  wire  mem_195_3_W0_clk;
  wire [7:0] mem_195_3_W0_data;
  wire  mem_195_3_W0_en;
  wire  mem_195_3_W0_mask;
  wire [25:0] mem_195_4_R0_addr;
  wire  mem_195_4_R0_clk;
  wire [7:0] mem_195_4_R0_data;
  wire  mem_195_4_R0_en;
  wire [25:0] mem_195_4_W0_addr;
  wire  mem_195_4_W0_clk;
  wire [7:0] mem_195_4_W0_data;
  wire  mem_195_4_W0_en;
  wire  mem_195_4_W0_mask;
  wire [25:0] mem_195_5_R0_addr;
  wire  mem_195_5_R0_clk;
  wire [7:0] mem_195_5_R0_data;
  wire  mem_195_5_R0_en;
  wire [25:0] mem_195_5_W0_addr;
  wire  mem_195_5_W0_clk;
  wire [7:0] mem_195_5_W0_data;
  wire  mem_195_5_W0_en;
  wire  mem_195_5_W0_mask;
  wire [25:0] mem_195_6_R0_addr;
  wire  mem_195_6_R0_clk;
  wire [7:0] mem_195_6_R0_data;
  wire  mem_195_6_R0_en;
  wire [25:0] mem_195_6_W0_addr;
  wire  mem_195_6_W0_clk;
  wire [7:0] mem_195_6_W0_data;
  wire  mem_195_6_W0_en;
  wire  mem_195_6_W0_mask;
  wire [25:0] mem_195_7_R0_addr;
  wire  mem_195_7_R0_clk;
  wire [7:0] mem_195_7_R0_data;
  wire  mem_195_7_R0_en;
  wire [25:0] mem_195_7_W0_addr;
  wire  mem_195_7_W0_clk;
  wire [7:0] mem_195_7_W0_data;
  wire  mem_195_7_W0_en;
  wire  mem_195_7_W0_mask;
  wire [25:0] mem_196_0_R0_addr;
  wire  mem_196_0_R0_clk;
  wire [7:0] mem_196_0_R0_data;
  wire  mem_196_0_R0_en;
  wire [25:0] mem_196_0_W0_addr;
  wire  mem_196_0_W0_clk;
  wire [7:0] mem_196_0_W0_data;
  wire  mem_196_0_W0_en;
  wire  mem_196_0_W0_mask;
  wire [25:0] mem_196_1_R0_addr;
  wire  mem_196_1_R0_clk;
  wire [7:0] mem_196_1_R0_data;
  wire  mem_196_1_R0_en;
  wire [25:0] mem_196_1_W0_addr;
  wire  mem_196_1_W0_clk;
  wire [7:0] mem_196_1_W0_data;
  wire  mem_196_1_W0_en;
  wire  mem_196_1_W0_mask;
  wire [25:0] mem_196_2_R0_addr;
  wire  mem_196_2_R0_clk;
  wire [7:0] mem_196_2_R0_data;
  wire  mem_196_2_R0_en;
  wire [25:0] mem_196_2_W0_addr;
  wire  mem_196_2_W0_clk;
  wire [7:0] mem_196_2_W0_data;
  wire  mem_196_2_W0_en;
  wire  mem_196_2_W0_mask;
  wire [25:0] mem_196_3_R0_addr;
  wire  mem_196_3_R0_clk;
  wire [7:0] mem_196_3_R0_data;
  wire  mem_196_3_R0_en;
  wire [25:0] mem_196_3_W0_addr;
  wire  mem_196_3_W0_clk;
  wire [7:0] mem_196_3_W0_data;
  wire  mem_196_3_W0_en;
  wire  mem_196_3_W0_mask;
  wire [25:0] mem_196_4_R0_addr;
  wire  mem_196_4_R0_clk;
  wire [7:0] mem_196_4_R0_data;
  wire  mem_196_4_R0_en;
  wire [25:0] mem_196_4_W0_addr;
  wire  mem_196_4_W0_clk;
  wire [7:0] mem_196_4_W0_data;
  wire  mem_196_4_W0_en;
  wire  mem_196_4_W0_mask;
  wire [25:0] mem_196_5_R0_addr;
  wire  mem_196_5_R0_clk;
  wire [7:0] mem_196_5_R0_data;
  wire  mem_196_5_R0_en;
  wire [25:0] mem_196_5_W0_addr;
  wire  mem_196_5_W0_clk;
  wire [7:0] mem_196_5_W0_data;
  wire  mem_196_5_W0_en;
  wire  mem_196_5_W0_mask;
  wire [25:0] mem_196_6_R0_addr;
  wire  mem_196_6_R0_clk;
  wire [7:0] mem_196_6_R0_data;
  wire  mem_196_6_R0_en;
  wire [25:0] mem_196_6_W0_addr;
  wire  mem_196_6_W0_clk;
  wire [7:0] mem_196_6_W0_data;
  wire  mem_196_6_W0_en;
  wire  mem_196_6_W0_mask;
  wire [25:0] mem_196_7_R0_addr;
  wire  mem_196_7_R0_clk;
  wire [7:0] mem_196_7_R0_data;
  wire  mem_196_7_R0_en;
  wire [25:0] mem_196_7_W0_addr;
  wire  mem_196_7_W0_clk;
  wire [7:0] mem_196_7_W0_data;
  wire  mem_196_7_W0_en;
  wire  mem_196_7_W0_mask;
  wire [25:0] mem_197_0_R0_addr;
  wire  mem_197_0_R0_clk;
  wire [7:0] mem_197_0_R0_data;
  wire  mem_197_0_R0_en;
  wire [25:0] mem_197_0_W0_addr;
  wire  mem_197_0_W0_clk;
  wire [7:0] mem_197_0_W0_data;
  wire  mem_197_0_W0_en;
  wire  mem_197_0_W0_mask;
  wire [25:0] mem_197_1_R0_addr;
  wire  mem_197_1_R0_clk;
  wire [7:0] mem_197_1_R0_data;
  wire  mem_197_1_R0_en;
  wire [25:0] mem_197_1_W0_addr;
  wire  mem_197_1_W0_clk;
  wire [7:0] mem_197_1_W0_data;
  wire  mem_197_1_W0_en;
  wire  mem_197_1_W0_mask;
  wire [25:0] mem_197_2_R0_addr;
  wire  mem_197_2_R0_clk;
  wire [7:0] mem_197_2_R0_data;
  wire  mem_197_2_R0_en;
  wire [25:0] mem_197_2_W0_addr;
  wire  mem_197_2_W0_clk;
  wire [7:0] mem_197_2_W0_data;
  wire  mem_197_2_W0_en;
  wire  mem_197_2_W0_mask;
  wire [25:0] mem_197_3_R0_addr;
  wire  mem_197_3_R0_clk;
  wire [7:0] mem_197_3_R0_data;
  wire  mem_197_3_R0_en;
  wire [25:0] mem_197_3_W0_addr;
  wire  mem_197_3_W0_clk;
  wire [7:0] mem_197_3_W0_data;
  wire  mem_197_3_W0_en;
  wire  mem_197_3_W0_mask;
  wire [25:0] mem_197_4_R0_addr;
  wire  mem_197_4_R0_clk;
  wire [7:0] mem_197_4_R0_data;
  wire  mem_197_4_R0_en;
  wire [25:0] mem_197_4_W0_addr;
  wire  mem_197_4_W0_clk;
  wire [7:0] mem_197_4_W0_data;
  wire  mem_197_4_W0_en;
  wire  mem_197_4_W0_mask;
  wire [25:0] mem_197_5_R0_addr;
  wire  mem_197_5_R0_clk;
  wire [7:0] mem_197_5_R0_data;
  wire  mem_197_5_R0_en;
  wire [25:0] mem_197_5_W0_addr;
  wire  mem_197_5_W0_clk;
  wire [7:0] mem_197_5_W0_data;
  wire  mem_197_5_W0_en;
  wire  mem_197_5_W0_mask;
  wire [25:0] mem_197_6_R0_addr;
  wire  mem_197_6_R0_clk;
  wire [7:0] mem_197_6_R0_data;
  wire  mem_197_6_R0_en;
  wire [25:0] mem_197_6_W0_addr;
  wire  mem_197_6_W0_clk;
  wire [7:0] mem_197_6_W0_data;
  wire  mem_197_6_W0_en;
  wire  mem_197_6_W0_mask;
  wire [25:0] mem_197_7_R0_addr;
  wire  mem_197_7_R0_clk;
  wire [7:0] mem_197_7_R0_data;
  wire  mem_197_7_R0_en;
  wire [25:0] mem_197_7_W0_addr;
  wire  mem_197_7_W0_clk;
  wire [7:0] mem_197_7_W0_data;
  wire  mem_197_7_W0_en;
  wire  mem_197_7_W0_mask;
  wire [25:0] mem_198_0_R0_addr;
  wire  mem_198_0_R0_clk;
  wire [7:0] mem_198_0_R0_data;
  wire  mem_198_0_R0_en;
  wire [25:0] mem_198_0_W0_addr;
  wire  mem_198_0_W0_clk;
  wire [7:0] mem_198_0_W0_data;
  wire  mem_198_0_W0_en;
  wire  mem_198_0_W0_mask;
  wire [25:0] mem_198_1_R0_addr;
  wire  mem_198_1_R0_clk;
  wire [7:0] mem_198_1_R0_data;
  wire  mem_198_1_R0_en;
  wire [25:0] mem_198_1_W0_addr;
  wire  mem_198_1_W0_clk;
  wire [7:0] mem_198_1_W0_data;
  wire  mem_198_1_W0_en;
  wire  mem_198_1_W0_mask;
  wire [25:0] mem_198_2_R0_addr;
  wire  mem_198_2_R0_clk;
  wire [7:0] mem_198_2_R0_data;
  wire  mem_198_2_R0_en;
  wire [25:0] mem_198_2_W0_addr;
  wire  mem_198_2_W0_clk;
  wire [7:0] mem_198_2_W0_data;
  wire  mem_198_2_W0_en;
  wire  mem_198_2_W0_mask;
  wire [25:0] mem_198_3_R0_addr;
  wire  mem_198_3_R0_clk;
  wire [7:0] mem_198_3_R0_data;
  wire  mem_198_3_R0_en;
  wire [25:0] mem_198_3_W0_addr;
  wire  mem_198_3_W0_clk;
  wire [7:0] mem_198_3_W0_data;
  wire  mem_198_3_W0_en;
  wire  mem_198_3_W0_mask;
  wire [25:0] mem_198_4_R0_addr;
  wire  mem_198_4_R0_clk;
  wire [7:0] mem_198_4_R0_data;
  wire  mem_198_4_R0_en;
  wire [25:0] mem_198_4_W0_addr;
  wire  mem_198_4_W0_clk;
  wire [7:0] mem_198_4_W0_data;
  wire  mem_198_4_W0_en;
  wire  mem_198_4_W0_mask;
  wire [25:0] mem_198_5_R0_addr;
  wire  mem_198_5_R0_clk;
  wire [7:0] mem_198_5_R0_data;
  wire  mem_198_5_R0_en;
  wire [25:0] mem_198_5_W0_addr;
  wire  mem_198_5_W0_clk;
  wire [7:0] mem_198_5_W0_data;
  wire  mem_198_5_W0_en;
  wire  mem_198_5_W0_mask;
  wire [25:0] mem_198_6_R0_addr;
  wire  mem_198_6_R0_clk;
  wire [7:0] mem_198_6_R0_data;
  wire  mem_198_6_R0_en;
  wire [25:0] mem_198_6_W0_addr;
  wire  mem_198_6_W0_clk;
  wire [7:0] mem_198_6_W0_data;
  wire  mem_198_6_W0_en;
  wire  mem_198_6_W0_mask;
  wire [25:0] mem_198_7_R0_addr;
  wire  mem_198_7_R0_clk;
  wire [7:0] mem_198_7_R0_data;
  wire  mem_198_7_R0_en;
  wire [25:0] mem_198_7_W0_addr;
  wire  mem_198_7_W0_clk;
  wire [7:0] mem_198_7_W0_data;
  wire  mem_198_7_W0_en;
  wire  mem_198_7_W0_mask;
  wire [25:0] mem_199_0_R0_addr;
  wire  mem_199_0_R0_clk;
  wire [7:0] mem_199_0_R0_data;
  wire  mem_199_0_R0_en;
  wire [25:0] mem_199_0_W0_addr;
  wire  mem_199_0_W0_clk;
  wire [7:0] mem_199_0_W0_data;
  wire  mem_199_0_W0_en;
  wire  mem_199_0_W0_mask;
  wire [25:0] mem_199_1_R0_addr;
  wire  mem_199_1_R0_clk;
  wire [7:0] mem_199_1_R0_data;
  wire  mem_199_1_R0_en;
  wire [25:0] mem_199_1_W0_addr;
  wire  mem_199_1_W0_clk;
  wire [7:0] mem_199_1_W0_data;
  wire  mem_199_1_W0_en;
  wire  mem_199_1_W0_mask;
  wire [25:0] mem_199_2_R0_addr;
  wire  mem_199_2_R0_clk;
  wire [7:0] mem_199_2_R0_data;
  wire  mem_199_2_R0_en;
  wire [25:0] mem_199_2_W0_addr;
  wire  mem_199_2_W0_clk;
  wire [7:0] mem_199_2_W0_data;
  wire  mem_199_2_W0_en;
  wire  mem_199_2_W0_mask;
  wire [25:0] mem_199_3_R0_addr;
  wire  mem_199_3_R0_clk;
  wire [7:0] mem_199_3_R0_data;
  wire  mem_199_3_R0_en;
  wire [25:0] mem_199_3_W0_addr;
  wire  mem_199_3_W0_clk;
  wire [7:0] mem_199_3_W0_data;
  wire  mem_199_3_W0_en;
  wire  mem_199_3_W0_mask;
  wire [25:0] mem_199_4_R0_addr;
  wire  mem_199_4_R0_clk;
  wire [7:0] mem_199_4_R0_data;
  wire  mem_199_4_R0_en;
  wire [25:0] mem_199_4_W0_addr;
  wire  mem_199_4_W0_clk;
  wire [7:0] mem_199_4_W0_data;
  wire  mem_199_4_W0_en;
  wire  mem_199_4_W0_mask;
  wire [25:0] mem_199_5_R0_addr;
  wire  mem_199_5_R0_clk;
  wire [7:0] mem_199_5_R0_data;
  wire  mem_199_5_R0_en;
  wire [25:0] mem_199_5_W0_addr;
  wire  mem_199_5_W0_clk;
  wire [7:0] mem_199_5_W0_data;
  wire  mem_199_5_W0_en;
  wire  mem_199_5_W0_mask;
  wire [25:0] mem_199_6_R0_addr;
  wire  mem_199_6_R0_clk;
  wire [7:0] mem_199_6_R0_data;
  wire  mem_199_6_R0_en;
  wire [25:0] mem_199_6_W0_addr;
  wire  mem_199_6_W0_clk;
  wire [7:0] mem_199_6_W0_data;
  wire  mem_199_6_W0_en;
  wire  mem_199_6_W0_mask;
  wire [25:0] mem_199_7_R0_addr;
  wire  mem_199_7_R0_clk;
  wire [7:0] mem_199_7_R0_data;
  wire  mem_199_7_R0_en;
  wire [25:0] mem_199_7_W0_addr;
  wire  mem_199_7_W0_clk;
  wire [7:0] mem_199_7_W0_data;
  wire  mem_199_7_W0_en;
  wire  mem_199_7_W0_mask;
  wire [25:0] mem_200_0_R0_addr;
  wire  mem_200_0_R0_clk;
  wire [7:0] mem_200_0_R0_data;
  wire  mem_200_0_R0_en;
  wire [25:0] mem_200_0_W0_addr;
  wire  mem_200_0_W0_clk;
  wire [7:0] mem_200_0_W0_data;
  wire  mem_200_0_W0_en;
  wire  mem_200_0_W0_mask;
  wire [25:0] mem_200_1_R0_addr;
  wire  mem_200_1_R0_clk;
  wire [7:0] mem_200_1_R0_data;
  wire  mem_200_1_R0_en;
  wire [25:0] mem_200_1_W0_addr;
  wire  mem_200_1_W0_clk;
  wire [7:0] mem_200_1_W0_data;
  wire  mem_200_1_W0_en;
  wire  mem_200_1_W0_mask;
  wire [25:0] mem_200_2_R0_addr;
  wire  mem_200_2_R0_clk;
  wire [7:0] mem_200_2_R0_data;
  wire  mem_200_2_R0_en;
  wire [25:0] mem_200_2_W0_addr;
  wire  mem_200_2_W0_clk;
  wire [7:0] mem_200_2_W0_data;
  wire  mem_200_2_W0_en;
  wire  mem_200_2_W0_mask;
  wire [25:0] mem_200_3_R0_addr;
  wire  mem_200_3_R0_clk;
  wire [7:0] mem_200_3_R0_data;
  wire  mem_200_3_R0_en;
  wire [25:0] mem_200_3_W0_addr;
  wire  mem_200_3_W0_clk;
  wire [7:0] mem_200_3_W0_data;
  wire  mem_200_3_W0_en;
  wire  mem_200_3_W0_mask;
  wire [25:0] mem_200_4_R0_addr;
  wire  mem_200_4_R0_clk;
  wire [7:0] mem_200_4_R0_data;
  wire  mem_200_4_R0_en;
  wire [25:0] mem_200_4_W0_addr;
  wire  mem_200_4_W0_clk;
  wire [7:0] mem_200_4_W0_data;
  wire  mem_200_4_W0_en;
  wire  mem_200_4_W0_mask;
  wire [25:0] mem_200_5_R0_addr;
  wire  mem_200_5_R0_clk;
  wire [7:0] mem_200_5_R0_data;
  wire  mem_200_5_R0_en;
  wire [25:0] mem_200_5_W0_addr;
  wire  mem_200_5_W0_clk;
  wire [7:0] mem_200_5_W0_data;
  wire  mem_200_5_W0_en;
  wire  mem_200_5_W0_mask;
  wire [25:0] mem_200_6_R0_addr;
  wire  mem_200_6_R0_clk;
  wire [7:0] mem_200_6_R0_data;
  wire  mem_200_6_R0_en;
  wire [25:0] mem_200_6_W0_addr;
  wire  mem_200_6_W0_clk;
  wire [7:0] mem_200_6_W0_data;
  wire  mem_200_6_W0_en;
  wire  mem_200_6_W0_mask;
  wire [25:0] mem_200_7_R0_addr;
  wire  mem_200_7_R0_clk;
  wire [7:0] mem_200_7_R0_data;
  wire  mem_200_7_R0_en;
  wire [25:0] mem_200_7_W0_addr;
  wire  mem_200_7_W0_clk;
  wire [7:0] mem_200_7_W0_data;
  wire  mem_200_7_W0_en;
  wire  mem_200_7_W0_mask;
  wire [25:0] mem_201_0_R0_addr;
  wire  mem_201_0_R0_clk;
  wire [7:0] mem_201_0_R0_data;
  wire  mem_201_0_R0_en;
  wire [25:0] mem_201_0_W0_addr;
  wire  mem_201_0_W0_clk;
  wire [7:0] mem_201_0_W0_data;
  wire  mem_201_0_W0_en;
  wire  mem_201_0_W0_mask;
  wire [25:0] mem_201_1_R0_addr;
  wire  mem_201_1_R0_clk;
  wire [7:0] mem_201_1_R0_data;
  wire  mem_201_1_R0_en;
  wire [25:0] mem_201_1_W0_addr;
  wire  mem_201_1_W0_clk;
  wire [7:0] mem_201_1_W0_data;
  wire  mem_201_1_W0_en;
  wire  mem_201_1_W0_mask;
  wire [25:0] mem_201_2_R0_addr;
  wire  mem_201_2_R0_clk;
  wire [7:0] mem_201_2_R0_data;
  wire  mem_201_2_R0_en;
  wire [25:0] mem_201_2_W0_addr;
  wire  mem_201_2_W0_clk;
  wire [7:0] mem_201_2_W0_data;
  wire  mem_201_2_W0_en;
  wire  mem_201_2_W0_mask;
  wire [25:0] mem_201_3_R0_addr;
  wire  mem_201_3_R0_clk;
  wire [7:0] mem_201_3_R0_data;
  wire  mem_201_3_R0_en;
  wire [25:0] mem_201_3_W0_addr;
  wire  mem_201_3_W0_clk;
  wire [7:0] mem_201_3_W0_data;
  wire  mem_201_3_W0_en;
  wire  mem_201_3_W0_mask;
  wire [25:0] mem_201_4_R0_addr;
  wire  mem_201_4_R0_clk;
  wire [7:0] mem_201_4_R0_data;
  wire  mem_201_4_R0_en;
  wire [25:0] mem_201_4_W0_addr;
  wire  mem_201_4_W0_clk;
  wire [7:0] mem_201_4_W0_data;
  wire  mem_201_4_W0_en;
  wire  mem_201_4_W0_mask;
  wire [25:0] mem_201_5_R0_addr;
  wire  mem_201_5_R0_clk;
  wire [7:0] mem_201_5_R0_data;
  wire  mem_201_5_R0_en;
  wire [25:0] mem_201_5_W0_addr;
  wire  mem_201_5_W0_clk;
  wire [7:0] mem_201_5_W0_data;
  wire  mem_201_5_W0_en;
  wire  mem_201_5_W0_mask;
  wire [25:0] mem_201_6_R0_addr;
  wire  mem_201_6_R0_clk;
  wire [7:0] mem_201_6_R0_data;
  wire  mem_201_6_R0_en;
  wire [25:0] mem_201_6_W0_addr;
  wire  mem_201_6_W0_clk;
  wire [7:0] mem_201_6_W0_data;
  wire  mem_201_6_W0_en;
  wire  mem_201_6_W0_mask;
  wire [25:0] mem_201_7_R0_addr;
  wire  mem_201_7_R0_clk;
  wire [7:0] mem_201_7_R0_data;
  wire  mem_201_7_R0_en;
  wire [25:0] mem_201_7_W0_addr;
  wire  mem_201_7_W0_clk;
  wire [7:0] mem_201_7_W0_data;
  wire  mem_201_7_W0_en;
  wire  mem_201_7_W0_mask;
  wire [25:0] mem_202_0_R0_addr;
  wire  mem_202_0_R0_clk;
  wire [7:0] mem_202_0_R0_data;
  wire  mem_202_0_R0_en;
  wire [25:0] mem_202_0_W0_addr;
  wire  mem_202_0_W0_clk;
  wire [7:0] mem_202_0_W0_data;
  wire  mem_202_0_W0_en;
  wire  mem_202_0_W0_mask;
  wire [25:0] mem_202_1_R0_addr;
  wire  mem_202_1_R0_clk;
  wire [7:0] mem_202_1_R0_data;
  wire  mem_202_1_R0_en;
  wire [25:0] mem_202_1_W0_addr;
  wire  mem_202_1_W0_clk;
  wire [7:0] mem_202_1_W0_data;
  wire  mem_202_1_W0_en;
  wire  mem_202_1_W0_mask;
  wire [25:0] mem_202_2_R0_addr;
  wire  mem_202_2_R0_clk;
  wire [7:0] mem_202_2_R0_data;
  wire  mem_202_2_R0_en;
  wire [25:0] mem_202_2_W0_addr;
  wire  mem_202_2_W0_clk;
  wire [7:0] mem_202_2_W0_data;
  wire  mem_202_2_W0_en;
  wire  mem_202_2_W0_mask;
  wire [25:0] mem_202_3_R0_addr;
  wire  mem_202_3_R0_clk;
  wire [7:0] mem_202_3_R0_data;
  wire  mem_202_3_R0_en;
  wire [25:0] mem_202_3_W0_addr;
  wire  mem_202_3_W0_clk;
  wire [7:0] mem_202_3_W0_data;
  wire  mem_202_3_W0_en;
  wire  mem_202_3_W0_mask;
  wire [25:0] mem_202_4_R0_addr;
  wire  mem_202_4_R0_clk;
  wire [7:0] mem_202_4_R0_data;
  wire  mem_202_4_R0_en;
  wire [25:0] mem_202_4_W0_addr;
  wire  mem_202_4_W0_clk;
  wire [7:0] mem_202_4_W0_data;
  wire  mem_202_4_W0_en;
  wire  mem_202_4_W0_mask;
  wire [25:0] mem_202_5_R0_addr;
  wire  mem_202_5_R0_clk;
  wire [7:0] mem_202_5_R0_data;
  wire  mem_202_5_R0_en;
  wire [25:0] mem_202_5_W0_addr;
  wire  mem_202_5_W0_clk;
  wire [7:0] mem_202_5_W0_data;
  wire  mem_202_5_W0_en;
  wire  mem_202_5_W0_mask;
  wire [25:0] mem_202_6_R0_addr;
  wire  mem_202_6_R0_clk;
  wire [7:0] mem_202_6_R0_data;
  wire  mem_202_6_R0_en;
  wire [25:0] mem_202_6_W0_addr;
  wire  mem_202_6_W0_clk;
  wire [7:0] mem_202_6_W0_data;
  wire  mem_202_6_W0_en;
  wire  mem_202_6_W0_mask;
  wire [25:0] mem_202_7_R0_addr;
  wire  mem_202_7_R0_clk;
  wire [7:0] mem_202_7_R0_data;
  wire  mem_202_7_R0_en;
  wire [25:0] mem_202_7_W0_addr;
  wire  mem_202_7_W0_clk;
  wire [7:0] mem_202_7_W0_data;
  wire  mem_202_7_W0_en;
  wire  mem_202_7_W0_mask;
  wire [25:0] mem_203_0_R0_addr;
  wire  mem_203_0_R0_clk;
  wire [7:0] mem_203_0_R0_data;
  wire  mem_203_0_R0_en;
  wire [25:0] mem_203_0_W0_addr;
  wire  mem_203_0_W0_clk;
  wire [7:0] mem_203_0_W0_data;
  wire  mem_203_0_W0_en;
  wire  mem_203_0_W0_mask;
  wire [25:0] mem_203_1_R0_addr;
  wire  mem_203_1_R0_clk;
  wire [7:0] mem_203_1_R0_data;
  wire  mem_203_1_R0_en;
  wire [25:0] mem_203_1_W0_addr;
  wire  mem_203_1_W0_clk;
  wire [7:0] mem_203_1_W0_data;
  wire  mem_203_1_W0_en;
  wire  mem_203_1_W0_mask;
  wire [25:0] mem_203_2_R0_addr;
  wire  mem_203_2_R0_clk;
  wire [7:0] mem_203_2_R0_data;
  wire  mem_203_2_R0_en;
  wire [25:0] mem_203_2_W0_addr;
  wire  mem_203_2_W0_clk;
  wire [7:0] mem_203_2_W0_data;
  wire  mem_203_2_W0_en;
  wire  mem_203_2_W0_mask;
  wire [25:0] mem_203_3_R0_addr;
  wire  mem_203_3_R0_clk;
  wire [7:0] mem_203_3_R0_data;
  wire  mem_203_3_R0_en;
  wire [25:0] mem_203_3_W0_addr;
  wire  mem_203_3_W0_clk;
  wire [7:0] mem_203_3_W0_data;
  wire  mem_203_3_W0_en;
  wire  mem_203_3_W0_mask;
  wire [25:0] mem_203_4_R0_addr;
  wire  mem_203_4_R0_clk;
  wire [7:0] mem_203_4_R0_data;
  wire  mem_203_4_R0_en;
  wire [25:0] mem_203_4_W0_addr;
  wire  mem_203_4_W0_clk;
  wire [7:0] mem_203_4_W0_data;
  wire  mem_203_4_W0_en;
  wire  mem_203_4_W0_mask;
  wire [25:0] mem_203_5_R0_addr;
  wire  mem_203_5_R0_clk;
  wire [7:0] mem_203_5_R0_data;
  wire  mem_203_5_R0_en;
  wire [25:0] mem_203_5_W0_addr;
  wire  mem_203_5_W0_clk;
  wire [7:0] mem_203_5_W0_data;
  wire  mem_203_5_W0_en;
  wire  mem_203_5_W0_mask;
  wire [25:0] mem_203_6_R0_addr;
  wire  mem_203_6_R0_clk;
  wire [7:0] mem_203_6_R0_data;
  wire  mem_203_6_R0_en;
  wire [25:0] mem_203_6_W0_addr;
  wire  mem_203_6_W0_clk;
  wire [7:0] mem_203_6_W0_data;
  wire  mem_203_6_W0_en;
  wire  mem_203_6_W0_mask;
  wire [25:0] mem_203_7_R0_addr;
  wire  mem_203_7_R0_clk;
  wire [7:0] mem_203_7_R0_data;
  wire  mem_203_7_R0_en;
  wire [25:0] mem_203_7_W0_addr;
  wire  mem_203_7_W0_clk;
  wire [7:0] mem_203_7_W0_data;
  wire  mem_203_7_W0_en;
  wire  mem_203_7_W0_mask;
  wire [25:0] mem_204_0_R0_addr;
  wire  mem_204_0_R0_clk;
  wire [7:0] mem_204_0_R0_data;
  wire  mem_204_0_R0_en;
  wire [25:0] mem_204_0_W0_addr;
  wire  mem_204_0_W0_clk;
  wire [7:0] mem_204_0_W0_data;
  wire  mem_204_0_W0_en;
  wire  mem_204_0_W0_mask;
  wire [25:0] mem_204_1_R0_addr;
  wire  mem_204_1_R0_clk;
  wire [7:0] mem_204_1_R0_data;
  wire  mem_204_1_R0_en;
  wire [25:0] mem_204_1_W0_addr;
  wire  mem_204_1_W0_clk;
  wire [7:0] mem_204_1_W0_data;
  wire  mem_204_1_W0_en;
  wire  mem_204_1_W0_mask;
  wire [25:0] mem_204_2_R0_addr;
  wire  mem_204_2_R0_clk;
  wire [7:0] mem_204_2_R0_data;
  wire  mem_204_2_R0_en;
  wire [25:0] mem_204_2_W0_addr;
  wire  mem_204_2_W0_clk;
  wire [7:0] mem_204_2_W0_data;
  wire  mem_204_2_W0_en;
  wire  mem_204_2_W0_mask;
  wire [25:0] mem_204_3_R0_addr;
  wire  mem_204_3_R0_clk;
  wire [7:0] mem_204_3_R0_data;
  wire  mem_204_3_R0_en;
  wire [25:0] mem_204_3_W0_addr;
  wire  mem_204_3_W0_clk;
  wire [7:0] mem_204_3_W0_data;
  wire  mem_204_3_W0_en;
  wire  mem_204_3_W0_mask;
  wire [25:0] mem_204_4_R0_addr;
  wire  mem_204_4_R0_clk;
  wire [7:0] mem_204_4_R0_data;
  wire  mem_204_4_R0_en;
  wire [25:0] mem_204_4_W0_addr;
  wire  mem_204_4_W0_clk;
  wire [7:0] mem_204_4_W0_data;
  wire  mem_204_4_W0_en;
  wire  mem_204_4_W0_mask;
  wire [25:0] mem_204_5_R0_addr;
  wire  mem_204_5_R0_clk;
  wire [7:0] mem_204_5_R0_data;
  wire  mem_204_5_R0_en;
  wire [25:0] mem_204_5_W0_addr;
  wire  mem_204_5_W0_clk;
  wire [7:0] mem_204_5_W0_data;
  wire  mem_204_5_W0_en;
  wire  mem_204_5_W0_mask;
  wire [25:0] mem_204_6_R0_addr;
  wire  mem_204_6_R0_clk;
  wire [7:0] mem_204_6_R0_data;
  wire  mem_204_6_R0_en;
  wire [25:0] mem_204_6_W0_addr;
  wire  mem_204_6_W0_clk;
  wire [7:0] mem_204_6_W0_data;
  wire  mem_204_6_W0_en;
  wire  mem_204_6_W0_mask;
  wire [25:0] mem_204_7_R0_addr;
  wire  mem_204_7_R0_clk;
  wire [7:0] mem_204_7_R0_data;
  wire  mem_204_7_R0_en;
  wire [25:0] mem_204_7_W0_addr;
  wire  mem_204_7_W0_clk;
  wire [7:0] mem_204_7_W0_data;
  wire  mem_204_7_W0_en;
  wire  mem_204_7_W0_mask;
  wire [25:0] mem_205_0_R0_addr;
  wire  mem_205_0_R0_clk;
  wire [7:0] mem_205_0_R0_data;
  wire  mem_205_0_R0_en;
  wire [25:0] mem_205_0_W0_addr;
  wire  mem_205_0_W0_clk;
  wire [7:0] mem_205_0_W0_data;
  wire  mem_205_0_W0_en;
  wire  mem_205_0_W0_mask;
  wire [25:0] mem_205_1_R0_addr;
  wire  mem_205_1_R0_clk;
  wire [7:0] mem_205_1_R0_data;
  wire  mem_205_1_R0_en;
  wire [25:0] mem_205_1_W0_addr;
  wire  mem_205_1_W0_clk;
  wire [7:0] mem_205_1_W0_data;
  wire  mem_205_1_W0_en;
  wire  mem_205_1_W0_mask;
  wire [25:0] mem_205_2_R0_addr;
  wire  mem_205_2_R0_clk;
  wire [7:0] mem_205_2_R0_data;
  wire  mem_205_2_R0_en;
  wire [25:0] mem_205_2_W0_addr;
  wire  mem_205_2_W0_clk;
  wire [7:0] mem_205_2_W0_data;
  wire  mem_205_2_W0_en;
  wire  mem_205_2_W0_mask;
  wire [25:0] mem_205_3_R0_addr;
  wire  mem_205_3_R0_clk;
  wire [7:0] mem_205_3_R0_data;
  wire  mem_205_3_R0_en;
  wire [25:0] mem_205_3_W0_addr;
  wire  mem_205_3_W0_clk;
  wire [7:0] mem_205_3_W0_data;
  wire  mem_205_3_W0_en;
  wire  mem_205_3_W0_mask;
  wire [25:0] mem_205_4_R0_addr;
  wire  mem_205_4_R0_clk;
  wire [7:0] mem_205_4_R0_data;
  wire  mem_205_4_R0_en;
  wire [25:0] mem_205_4_W0_addr;
  wire  mem_205_4_W0_clk;
  wire [7:0] mem_205_4_W0_data;
  wire  mem_205_4_W0_en;
  wire  mem_205_4_W0_mask;
  wire [25:0] mem_205_5_R0_addr;
  wire  mem_205_5_R0_clk;
  wire [7:0] mem_205_5_R0_data;
  wire  mem_205_5_R0_en;
  wire [25:0] mem_205_5_W0_addr;
  wire  mem_205_5_W0_clk;
  wire [7:0] mem_205_5_W0_data;
  wire  mem_205_5_W0_en;
  wire  mem_205_5_W0_mask;
  wire [25:0] mem_205_6_R0_addr;
  wire  mem_205_6_R0_clk;
  wire [7:0] mem_205_6_R0_data;
  wire  mem_205_6_R0_en;
  wire [25:0] mem_205_6_W0_addr;
  wire  mem_205_6_W0_clk;
  wire [7:0] mem_205_6_W0_data;
  wire  mem_205_6_W0_en;
  wire  mem_205_6_W0_mask;
  wire [25:0] mem_205_7_R0_addr;
  wire  mem_205_7_R0_clk;
  wire [7:0] mem_205_7_R0_data;
  wire  mem_205_7_R0_en;
  wire [25:0] mem_205_7_W0_addr;
  wire  mem_205_7_W0_clk;
  wire [7:0] mem_205_7_W0_data;
  wire  mem_205_7_W0_en;
  wire  mem_205_7_W0_mask;
  wire [25:0] mem_206_0_R0_addr;
  wire  mem_206_0_R0_clk;
  wire [7:0] mem_206_0_R0_data;
  wire  mem_206_0_R0_en;
  wire [25:0] mem_206_0_W0_addr;
  wire  mem_206_0_W0_clk;
  wire [7:0] mem_206_0_W0_data;
  wire  mem_206_0_W0_en;
  wire  mem_206_0_W0_mask;
  wire [25:0] mem_206_1_R0_addr;
  wire  mem_206_1_R0_clk;
  wire [7:0] mem_206_1_R0_data;
  wire  mem_206_1_R0_en;
  wire [25:0] mem_206_1_W0_addr;
  wire  mem_206_1_W0_clk;
  wire [7:0] mem_206_1_W0_data;
  wire  mem_206_1_W0_en;
  wire  mem_206_1_W0_mask;
  wire [25:0] mem_206_2_R0_addr;
  wire  mem_206_2_R0_clk;
  wire [7:0] mem_206_2_R0_data;
  wire  mem_206_2_R0_en;
  wire [25:0] mem_206_2_W0_addr;
  wire  mem_206_2_W0_clk;
  wire [7:0] mem_206_2_W0_data;
  wire  mem_206_2_W0_en;
  wire  mem_206_2_W0_mask;
  wire [25:0] mem_206_3_R0_addr;
  wire  mem_206_3_R0_clk;
  wire [7:0] mem_206_3_R0_data;
  wire  mem_206_3_R0_en;
  wire [25:0] mem_206_3_W0_addr;
  wire  mem_206_3_W0_clk;
  wire [7:0] mem_206_3_W0_data;
  wire  mem_206_3_W0_en;
  wire  mem_206_3_W0_mask;
  wire [25:0] mem_206_4_R0_addr;
  wire  mem_206_4_R0_clk;
  wire [7:0] mem_206_4_R0_data;
  wire  mem_206_4_R0_en;
  wire [25:0] mem_206_4_W0_addr;
  wire  mem_206_4_W0_clk;
  wire [7:0] mem_206_4_W0_data;
  wire  mem_206_4_W0_en;
  wire  mem_206_4_W0_mask;
  wire [25:0] mem_206_5_R0_addr;
  wire  mem_206_5_R0_clk;
  wire [7:0] mem_206_5_R0_data;
  wire  mem_206_5_R0_en;
  wire [25:0] mem_206_5_W0_addr;
  wire  mem_206_5_W0_clk;
  wire [7:0] mem_206_5_W0_data;
  wire  mem_206_5_W0_en;
  wire  mem_206_5_W0_mask;
  wire [25:0] mem_206_6_R0_addr;
  wire  mem_206_6_R0_clk;
  wire [7:0] mem_206_6_R0_data;
  wire  mem_206_6_R0_en;
  wire [25:0] mem_206_6_W0_addr;
  wire  mem_206_6_W0_clk;
  wire [7:0] mem_206_6_W0_data;
  wire  mem_206_6_W0_en;
  wire  mem_206_6_W0_mask;
  wire [25:0] mem_206_7_R0_addr;
  wire  mem_206_7_R0_clk;
  wire [7:0] mem_206_7_R0_data;
  wire  mem_206_7_R0_en;
  wire [25:0] mem_206_7_W0_addr;
  wire  mem_206_7_W0_clk;
  wire [7:0] mem_206_7_W0_data;
  wire  mem_206_7_W0_en;
  wire  mem_206_7_W0_mask;
  wire [25:0] mem_207_0_R0_addr;
  wire  mem_207_0_R0_clk;
  wire [7:0] mem_207_0_R0_data;
  wire  mem_207_0_R0_en;
  wire [25:0] mem_207_0_W0_addr;
  wire  mem_207_0_W0_clk;
  wire [7:0] mem_207_0_W0_data;
  wire  mem_207_0_W0_en;
  wire  mem_207_0_W0_mask;
  wire [25:0] mem_207_1_R0_addr;
  wire  mem_207_1_R0_clk;
  wire [7:0] mem_207_1_R0_data;
  wire  mem_207_1_R0_en;
  wire [25:0] mem_207_1_W0_addr;
  wire  mem_207_1_W0_clk;
  wire [7:0] mem_207_1_W0_data;
  wire  mem_207_1_W0_en;
  wire  mem_207_1_W0_mask;
  wire [25:0] mem_207_2_R0_addr;
  wire  mem_207_2_R0_clk;
  wire [7:0] mem_207_2_R0_data;
  wire  mem_207_2_R0_en;
  wire [25:0] mem_207_2_W0_addr;
  wire  mem_207_2_W0_clk;
  wire [7:0] mem_207_2_W0_data;
  wire  mem_207_2_W0_en;
  wire  mem_207_2_W0_mask;
  wire [25:0] mem_207_3_R0_addr;
  wire  mem_207_3_R0_clk;
  wire [7:0] mem_207_3_R0_data;
  wire  mem_207_3_R0_en;
  wire [25:0] mem_207_3_W0_addr;
  wire  mem_207_3_W0_clk;
  wire [7:0] mem_207_3_W0_data;
  wire  mem_207_3_W0_en;
  wire  mem_207_3_W0_mask;
  wire [25:0] mem_207_4_R0_addr;
  wire  mem_207_4_R0_clk;
  wire [7:0] mem_207_4_R0_data;
  wire  mem_207_4_R0_en;
  wire [25:0] mem_207_4_W0_addr;
  wire  mem_207_4_W0_clk;
  wire [7:0] mem_207_4_W0_data;
  wire  mem_207_4_W0_en;
  wire  mem_207_4_W0_mask;
  wire [25:0] mem_207_5_R0_addr;
  wire  mem_207_5_R0_clk;
  wire [7:0] mem_207_5_R0_data;
  wire  mem_207_5_R0_en;
  wire [25:0] mem_207_5_W0_addr;
  wire  mem_207_5_W0_clk;
  wire [7:0] mem_207_5_W0_data;
  wire  mem_207_5_W0_en;
  wire  mem_207_5_W0_mask;
  wire [25:0] mem_207_6_R0_addr;
  wire  mem_207_6_R0_clk;
  wire [7:0] mem_207_6_R0_data;
  wire  mem_207_6_R0_en;
  wire [25:0] mem_207_6_W0_addr;
  wire  mem_207_6_W0_clk;
  wire [7:0] mem_207_6_W0_data;
  wire  mem_207_6_W0_en;
  wire  mem_207_6_W0_mask;
  wire [25:0] mem_207_7_R0_addr;
  wire  mem_207_7_R0_clk;
  wire [7:0] mem_207_7_R0_data;
  wire  mem_207_7_R0_en;
  wire [25:0] mem_207_7_W0_addr;
  wire  mem_207_7_W0_clk;
  wire [7:0] mem_207_7_W0_data;
  wire  mem_207_7_W0_en;
  wire  mem_207_7_W0_mask;
  wire [25:0] mem_208_0_R0_addr;
  wire  mem_208_0_R0_clk;
  wire [7:0] mem_208_0_R0_data;
  wire  mem_208_0_R0_en;
  wire [25:0] mem_208_0_W0_addr;
  wire  mem_208_0_W0_clk;
  wire [7:0] mem_208_0_W0_data;
  wire  mem_208_0_W0_en;
  wire  mem_208_0_W0_mask;
  wire [25:0] mem_208_1_R0_addr;
  wire  mem_208_1_R0_clk;
  wire [7:0] mem_208_1_R0_data;
  wire  mem_208_1_R0_en;
  wire [25:0] mem_208_1_W0_addr;
  wire  mem_208_1_W0_clk;
  wire [7:0] mem_208_1_W0_data;
  wire  mem_208_1_W0_en;
  wire  mem_208_1_W0_mask;
  wire [25:0] mem_208_2_R0_addr;
  wire  mem_208_2_R0_clk;
  wire [7:0] mem_208_2_R0_data;
  wire  mem_208_2_R0_en;
  wire [25:0] mem_208_2_W0_addr;
  wire  mem_208_2_W0_clk;
  wire [7:0] mem_208_2_W0_data;
  wire  mem_208_2_W0_en;
  wire  mem_208_2_W0_mask;
  wire [25:0] mem_208_3_R0_addr;
  wire  mem_208_3_R0_clk;
  wire [7:0] mem_208_3_R0_data;
  wire  mem_208_3_R0_en;
  wire [25:0] mem_208_3_W0_addr;
  wire  mem_208_3_W0_clk;
  wire [7:0] mem_208_3_W0_data;
  wire  mem_208_3_W0_en;
  wire  mem_208_3_W0_mask;
  wire [25:0] mem_208_4_R0_addr;
  wire  mem_208_4_R0_clk;
  wire [7:0] mem_208_4_R0_data;
  wire  mem_208_4_R0_en;
  wire [25:0] mem_208_4_W0_addr;
  wire  mem_208_4_W0_clk;
  wire [7:0] mem_208_4_W0_data;
  wire  mem_208_4_W0_en;
  wire  mem_208_4_W0_mask;
  wire [25:0] mem_208_5_R0_addr;
  wire  mem_208_5_R0_clk;
  wire [7:0] mem_208_5_R0_data;
  wire  mem_208_5_R0_en;
  wire [25:0] mem_208_5_W0_addr;
  wire  mem_208_5_W0_clk;
  wire [7:0] mem_208_5_W0_data;
  wire  mem_208_5_W0_en;
  wire  mem_208_5_W0_mask;
  wire [25:0] mem_208_6_R0_addr;
  wire  mem_208_6_R0_clk;
  wire [7:0] mem_208_6_R0_data;
  wire  mem_208_6_R0_en;
  wire [25:0] mem_208_6_W0_addr;
  wire  mem_208_6_W0_clk;
  wire [7:0] mem_208_6_W0_data;
  wire  mem_208_6_W0_en;
  wire  mem_208_6_W0_mask;
  wire [25:0] mem_208_7_R0_addr;
  wire  mem_208_7_R0_clk;
  wire [7:0] mem_208_7_R0_data;
  wire  mem_208_7_R0_en;
  wire [25:0] mem_208_7_W0_addr;
  wire  mem_208_7_W0_clk;
  wire [7:0] mem_208_7_W0_data;
  wire  mem_208_7_W0_en;
  wire  mem_208_7_W0_mask;
  wire [25:0] mem_209_0_R0_addr;
  wire  mem_209_0_R0_clk;
  wire [7:0] mem_209_0_R0_data;
  wire  mem_209_0_R0_en;
  wire [25:0] mem_209_0_W0_addr;
  wire  mem_209_0_W0_clk;
  wire [7:0] mem_209_0_W0_data;
  wire  mem_209_0_W0_en;
  wire  mem_209_0_W0_mask;
  wire [25:0] mem_209_1_R0_addr;
  wire  mem_209_1_R0_clk;
  wire [7:0] mem_209_1_R0_data;
  wire  mem_209_1_R0_en;
  wire [25:0] mem_209_1_W0_addr;
  wire  mem_209_1_W0_clk;
  wire [7:0] mem_209_1_W0_data;
  wire  mem_209_1_W0_en;
  wire  mem_209_1_W0_mask;
  wire [25:0] mem_209_2_R0_addr;
  wire  mem_209_2_R0_clk;
  wire [7:0] mem_209_2_R0_data;
  wire  mem_209_2_R0_en;
  wire [25:0] mem_209_2_W0_addr;
  wire  mem_209_2_W0_clk;
  wire [7:0] mem_209_2_W0_data;
  wire  mem_209_2_W0_en;
  wire  mem_209_2_W0_mask;
  wire [25:0] mem_209_3_R0_addr;
  wire  mem_209_3_R0_clk;
  wire [7:0] mem_209_3_R0_data;
  wire  mem_209_3_R0_en;
  wire [25:0] mem_209_3_W0_addr;
  wire  mem_209_3_W0_clk;
  wire [7:0] mem_209_3_W0_data;
  wire  mem_209_3_W0_en;
  wire  mem_209_3_W0_mask;
  wire [25:0] mem_209_4_R0_addr;
  wire  mem_209_4_R0_clk;
  wire [7:0] mem_209_4_R0_data;
  wire  mem_209_4_R0_en;
  wire [25:0] mem_209_4_W0_addr;
  wire  mem_209_4_W0_clk;
  wire [7:0] mem_209_4_W0_data;
  wire  mem_209_4_W0_en;
  wire  mem_209_4_W0_mask;
  wire [25:0] mem_209_5_R0_addr;
  wire  mem_209_5_R0_clk;
  wire [7:0] mem_209_5_R0_data;
  wire  mem_209_5_R0_en;
  wire [25:0] mem_209_5_W0_addr;
  wire  mem_209_5_W0_clk;
  wire [7:0] mem_209_5_W0_data;
  wire  mem_209_5_W0_en;
  wire  mem_209_5_W0_mask;
  wire [25:0] mem_209_6_R0_addr;
  wire  mem_209_6_R0_clk;
  wire [7:0] mem_209_6_R0_data;
  wire  mem_209_6_R0_en;
  wire [25:0] mem_209_6_W0_addr;
  wire  mem_209_6_W0_clk;
  wire [7:0] mem_209_6_W0_data;
  wire  mem_209_6_W0_en;
  wire  mem_209_6_W0_mask;
  wire [25:0] mem_209_7_R0_addr;
  wire  mem_209_7_R0_clk;
  wire [7:0] mem_209_7_R0_data;
  wire  mem_209_7_R0_en;
  wire [25:0] mem_209_7_W0_addr;
  wire  mem_209_7_W0_clk;
  wire [7:0] mem_209_7_W0_data;
  wire  mem_209_7_W0_en;
  wire  mem_209_7_W0_mask;
  wire [25:0] mem_210_0_R0_addr;
  wire  mem_210_0_R0_clk;
  wire [7:0] mem_210_0_R0_data;
  wire  mem_210_0_R0_en;
  wire [25:0] mem_210_0_W0_addr;
  wire  mem_210_0_W0_clk;
  wire [7:0] mem_210_0_W0_data;
  wire  mem_210_0_W0_en;
  wire  mem_210_0_W0_mask;
  wire [25:0] mem_210_1_R0_addr;
  wire  mem_210_1_R0_clk;
  wire [7:0] mem_210_1_R0_data;
  wire  mem_210_1_R0_en;
  wire [25:0] mem_210_1_W0_addr;
  wire  mem_210_1_W0_clk;
  wire [7:0] mem_210_1_W0_data;
  wire  mem_210_1_W0_en;
  wire  mem_210_1_W0_mask;
  wire [25:0] mem_210_2_R0_addr;
  wire  mem_210_2_R0_clk;
  wire [7:0] mem_210_2_R0_data;
  wire  mem_210_2_R0_en;
  wire [25:0] mem_210_2_W0_addr;
  wire  mem_210_2_W0_clk;
  wire [7:0] mem_210_2_W0_data;
  wire  mem_210_2_W0_en;
  wire  mem_210_2_W0_mask;
  wire [25:0] mem_210_3_R0_addr;
  wire  mem_210_3_R0_clk;
  wire [7:0] mem_210_3_R0_data;
  wire  mem_210_3_R0_en;
  wire [25:0] mem_210_3_W0_addr;
  wire  mem_210_3_W0_clk;
  wire [7:0] mem_210_3_W0_data;
  wire  mem_210_3_W0_en;
  wire  mem_210_3_W0_mask;
  wire [25:0] mem_210_4_R0_addr;
  wire  mem_210_4_R0_clk;
  wire [7:0] mem_210_4_R0_data;
  wire  mem_210_4_R0_en;
  wire [25:0] mem_210_4_W0_addr;
  wire  mem_210_4_W0_clk;
  wire [7:0] mem_210_4_W0_data;
  wire  mem_210_4_W0_en;
  wire  mem_210_4_W0_mask;
  wire [25:0] mem_210_5_R0_addr;
  wire  mem_210_5_R0_clk;
  wire [7:0] mem_210_5_R0_data;
  wire  mem_210_5_R0_en;
  wire [25:0] mem_210_5_W0_addr;
  wire  mem_210_5_W0_clk;
  wire [7:0] mem_210_5_W0_data;
  wire  mem_210_5_W0_en;
  wire  mem_210_5_W0_mask;
  wire [25:0] mem_210_6_R0_addr;
  wire  mem_210_6_R0_clk;
  wire [7:0] mem_210_6_R0_data;
  wire  mem_210_6_R0_en;
  wire [25:0] mem_210_6_W0_addr;
  wire  mem_210_6_W0_clk;
  wire [7:0] mem_210_6_W0_data;
  wire  mem_210_6_W0_en;
  wire  mem_210_6_W0_mask;
  wire [25:0] mem_210_7_R0_addr;
  wire  mem_210_7_R0_clk;
  wire [7:0] mem_210_7_R0_data;
  wire  mem_210_7_R0_en;
  wire [25:0] mem_210_7_W0_addr;
  wire  mem_210_7_W0_clk;
  wire [7:0] mem_210_7_W0_data;
  wire  mem_210_7_W0_en;
  wire  mem_210_7_W0_mask;
  wire [25:0] mem_211_0_R0_addr;
  wire  mem_211_0_R0_clk;
  wire [7:0] mem_211_0_R0_data;
  wire  mem_211_0_R0_en;
  wire [25:0] mem_211_0_W0_addr;
  wire  mem_211_0_W0_clk;
  wire [7:0] mem_211_0_W0_data;
  wire  mem_211_0_W0_en;
  wire  mem_211_0_W0_mask;
  wire [25:0] mem_211_1_R0_addr;
  wire  mem_211_1_R0_clk;
  wire [7:0] mem_211_1_R0_data;
  wire  mem_211_1_R0_en;
  wire [25:0] mem_211_1_W0_addr;
  wire  mem_211_1_W0_clk;
  wire [7:0] mem_211_1_W0_data;
  wire  mem_211_1_W0_en;
  wire  mem_211_1_W0_mask;
  wire [25:0] mem_211_2_R0_addr;
  wire  mem_211_2_R0_clk;
  wire [7:0] mem_211_2_R0_data;
  wire  mem_211_2_R0_en;
  wire [25:0] mem_211_2_W0_addr;
  wire  mem_211_2_W0_clk;
  wire [7:0] mem_211_2_W0_data;
  wire  mem_211_2_W0_en;
  wire  mem_211_2_W0_mask;
  wire [25:0] mem_211_3_R0_addr;
  wire  mem_211_3_R0_clk;
  wire [7:0] mem_211_3_R0_data;
  wire  mem_211_3_R0_en;
  wire [25:0] mem_211_3_W0_addr;
  wire  mem_211_3_W0_clk;
  wire [7:0] mem_211_3_W0_data;
  wire  mem_211_3_W0_en;
  wire  mem_211_3_W0_mask;
  wire [25:0] mem_211_4_R0_addr;
  wire  mem_211_4_R0_clk;
  wire [7:0] mem_211_4_R0_data;
  wire  mem_211_4_R0_en;
  wire [25:0] mem_211_4_W0_addr;
  wire  mem_211_4_W0_clk;
  wire [7:0] mem_211_4_W0_data;
  wire  mem_211_4_W0_en;
  wire  mem_211_4_W0_mask;
  wire [25:0] mem_211_5_R0_addr;
  wire  mem_211_5_R0_clk;
  wire [7:0] mem_211_5_R0_data;
  wire  mem_211_5_R0_en;
  wire [25:0] mem_211_5_W0_addr;
  wire  mem_211_5_W0_clk;
  wire [7:0] mem_211_5_W0_data;
  wire  mem_211_5_W0_en;
  wire  mem_211_5_W0_mask;
  wire [25:0] mem_211_6_R0_addr;
  wire  mem_211_6_R0_clk;
  wire [7:0] mem_211_6_R0_data;
  wire  mem_211_6_R0_en;
  wire [25:0] mem_211_6_W0_addr;
  wire  mem_211_6_W0_clk;
  wire [7:0] mem_211_6_W0_data;
  wire  mem_211_6_W0_en;
  wire  mem_211_6_W0_mask;
  wire [25:0] mem_211_7_R0_addr;
  wire  mem_211_7_R0_clk;
  wire [7:0] mem_211_7_R0_data;
  wire  mem_211_7_R0_en;
  wire [25:0] mem_211_7_W0_addr;
  wire  mem_211_7_W0_clk;
  wire [7:0] mem_211_7_W0_data;
  wire  mem_211_7_W0_en;
  wire  mem_211_7_W0_mask;
  wire [25:0] mem_212_0_R0_addr;
  wire  mem_212_0_R0_clk;
  wire [7:0] mem_212_0_R0_data;
  wire  mem_212_0_R0_en;
  wire [25:0] mem_212_0_W0_addr;
  wire  mem_212_0_W0_clk;
  wire [7:0] mem_212_0_W0_data;
  wire  mem_212_0_W0_en;
  wire  mem_212_0_W0_mask;
  wire [25:0] mem_212_1_R0_addr;
  wire  mem_212_1_R0_clk;
  wire [7:0] mem_212_1_R0_data;
  wire  mem_212_1_R0_en;
  wire [25:0] mem_212_1_W0_addr;
  wire  mem_212_1_W0_clk;
  wire [7:0] mem_212_1_W0_data;
  wire  mem_212_1_W0_en;
  wire  mem_212_1_W0_mask;
  wire [25:0] mem_212_2_R0_addr;
  wire  mem_212_2_R0_clk;
  wire [7:0] mem_212_2_R0_data;
  wire  mem_212_2_R0_en;
  wire [25:0] mem_212_2_W0_addr;
  wire  mem_212_2_W0_clk;
  wire [7:0] mem_212_2_W0_data;
  wire  mem_212_2_W0_en;
  wire  mem_212_2_W0_mask;
  wire [25:0] mem_212_3_R0_addr;
  wire  mem_212_3_R0_clk;
  wire [7:0] mem_212_3_R0_data;
  wire  mem_212_3_R0_en;
  wire [25:0] mem_212_3_W0_addr;
  wire  mem_212_3_W0_clk;
  wire [7:0] mem_212_3_W0_data;
  wire  mem_212_3_W0_en;
  wire  mem_212_3_W0_mask;
  wire [25:0] mem_212_4_R0_addr;
  wire  mem_212_4_R0_clk;
  wire [7:0] mem_212_4_R0_data;
  wire  mem_212_4_R0_en;
  wire [25:0] mem_212_4_W0_addr;
  wire  mem_212_4_W0_clk;
  wire [7:0] mem_212_4_W0_data;
  wire  mem_212_4_W0_en;
  wire  mem_212_4_W0_mask;
  wire [25:0] mem_212_5_R0_addr;
  wire  mem_212_5_R0_clk;
  wire [7:0] mem_212_5_R0_data;
  wire  mem_212_5_R0_en;
  wire [25:0] mem_212_5_W0_addr;
  wire  mem_212_5_W0_clk;
  wire [7:0] mem_212_5_W0_data;
  wire  mem_212_5_W0_en;
  wire  mem_212_5_W0_mask;
  wire [25:0] mem_212_6_R0_addr;
  wire  mem_212_6_R0_clk;
  wire [7:0] mem_212_6_R0_data;
  wire  mem_212_6_R0_en;
  wire [25:0] mem_212_6_W0_addr;
  wire  mem_212_6_W0_clk;
  wire [7:0] mem_212_6_W0_data;
  wire  mem_212_6_W0_en;
  wire  mem_212_6_W0_mask;
  wire [25:0] mem_212_7_R0_addr;
  wire  mem_212_7_R0_clk;
  wire [7:0] mem_212_7_R0_data;
  wire  mem_212_7_R0_en;
  wire [25:0] mem_212_7_W0_addr;
  wire  mem_212_7_W0_clk;
  wire [7:0] mem_212_7_W0_data;
  wire  mem_212_7_W0_en;
  wire  mem_212_7_W0_mask;
  wire [25:0] mem_213_0_R0_addr;
  wire  mem_213_0_R0_clk;
  wire [7:0] mem_213_0_R0_data;
  wire  mem_213_0_R0_en;
  wire [25:0] mem_213_0_W0_addr;
  wire  mem_213_0_W0_clk;
  wire [7:0] mem_213_0_W0_data;
  wire  mem_213_0_W0_en;
  wire  mem_213_0_W0_mask;
  wire [25:0] mem_213_1_R0_addr;
  wire  mem_213_1_R0_clk;
  wire [7:0] mem_213_1_R0_data;
  wire  mem_213_1_R0_en;
  wire [25:0] mem_213_1_W0_addr;
  wire  mem_213_1_W0_clk;
  wire [7:0] mem_213_1_W0_data;
  wire  mem_213_1_W0_en;
  wire  mem_213_1_W0_mask;
  wire [25:0] mem_213_2_R0_addr;
  wire  mem_213_2_R0_clk;
  wire [7:0] mem_213_2_R0_data;
  wire  mem_213_2_R0_en;
  wire [25:0] mem_213_2_W0_addr;
  wire  mem_213_2_W0_clk;
  wire [7:0] mem_213_2_W0_data;
  wire  mem_213_2_W0_en;
  wire  mem_213_2_W0_mask;
  wire [25:0] mem_213_3_R0_addr;
  wire  mem_213_3_R0_clk;
  wire [7:0] mem_213_3_R0_data;
  wire  mem_213_3_R0_en;
  wire [25:0] mem_213_3_W0_addr;
  wire  mem_213_3_W0_clk;
  wire [7:0] mem_213_3_W0_data;
  wire  mem_213_3_W0_en;
  wire  mem_213_3_W0_mask;
  wire [25:0] mem_213_4_R0_addr;
  wire  mem_213_4_R0_clk;
  wire [7:0] mem_213_4_R0_data;
  wire  mem_213_4_R0_en;
  wire [25:0] mem_213_4_W0_addr;
  wire  mem_213_4_W0_clk;
  wire [7:0] mem_213_4_W0_data;
  wire  mem_213_4_W0_en;
  wire  mem_213_4_W0_mask;
  wire [25:0] mem_213_5_R0_addr;
  wire  mem_213_5_R0_clk;
  wire [7:0] mem_213_5_R0_data;
  wire  mem_213_5_R0_en;
  wire [25:0] mem_213_5_W0_addr;
  wire  mem_213_5_W0_clk;
  wire [7:0] mem_213_5_W0_data;
  wire  mem_213_5_W0_en;
  wire  mem_213_5_W0_mask;
  wire [25:0] mem_213_6_R0_addr;
  wire  mem_213_6_R0_clk;
  wire [7:0] mem_213_6_R0_data;
  wire  mem_213_6_R0_en;
  wire [25:0] mem_213_6_W0_addr;
  wire  mem_213_6_W0_clk;
  wire [7:0] mem_213_6_W0_data;
  wire  mem_213_6_W0_en;
  wire  mem_213_6_W0_mask;
  wire [25:0] mem_213_7_R0_addr;
  wire  mem_213_7_R0_clk;
  wire [7:0] mem_213_7_R0_data;
  wire  mem_213_7_R0_en;
  wire [25:0] mem_213_7_W0_addr;
  wire  mem_213_7_W0_clk;
  wire [7:0] mem_213_7_W0_data;
  wire  mem_213_7_W0_en;
  wire  mem_213_7_W0_mask;
  wire [25:0] mem_214_0_R0_addr;
  wire  mem_214_0_R0_clk;
  wire [7:0] mem_214_0_R0_data;
  wire  mem_214_0_R0_en;
  wire [25:0] mem_214_0_W0_addr;
  wire  mem_214_0_W0_clk;
  wire [7:0] mem_214_0_W0_data;
  wire  mem_214_0_W0_en;
  wire  mem_214_0_W0_mask;
  wire [25:0] mem_214_1_R0_addr;
  wire  mem_214_1_R0_clk;
  wire [7:0] mem_214_1_R0_data;
  wire  mem_214_1_R0_en;
  wire [25:0] mem_214_1_W0_addr;
  wire  mem_214_1_W0_clk;
  wire [7:0] mem_214_1_W0_data;
  wire  mem_214_1_W0_en;
  wire  mem_214_1_W0_mask;
  wire [25:0] mem_214_2_R0_addr;
  wire  mem_214_2_R0_clk;
  wire [7:0] mem_214_2_R0_data;
  wire  mem_214_2_R0_en;
  wire [25:0] mem_214_2_W0_addr;
  wire  mem_214_2_W0_clk;
  wire [7:0] mem_214_2_W0_data;
  wire  mem_214_2_W0_en;
  wire  mem_214_2_W0_mask;
  wire [25:0] mem_214_3_R0_addr;
  wire  mem_214_3_R0_clk;
  wire [7:0] mem_214_3_R0_data;
  wire  mem_214_3_R0_en;
  wire [25:0] mem_214_3_W0_addr;
  wire  mem_214_3_W0_clk;
  wire [7:0] mem_214_3_W0_data;
  wire  mem_214_3_W0_en;
  wire  mem_214_3_W0_mask;
  wire [25:0] mem_214_4_R0_addr;
  wire  mem_214_4_R0_clk;
  wire [7:0] mem_214_4_R0_data;
  wire  mem_214_4_R0_en;
  wire [25:0] mem_214_4_W0_addr;
  wire  mem_214_4_W0_clk;
  wire [7:0] mem_214_4_W0_data;
  wire  mem_214_4_W0_en;
  wire  mem_214_4_W0_mask;
  wire [25:0] mem_214_5_R0_addr;
  wire  mem_214_5_R0_clk;
  wire [7:0] mem_214_5_R0_data;
  wire  mem_214_5_R0_en;
  wire [25:0] mem_214_5_W0_addr;
  wire  mem_214_5_W0_clk;
  wire [7:0] mem_214_5_W0_data;
  wire  mem_214_5_W0_en;
  wire  mem_214_5_W0_mask;
  wire [25:0] mem_214_6_R0_addr;
  wire  mem_214_6_R0_clk;
  wire [7:0] mem_214_6_R0_data;
  wire  mem_214_6_R0_en;
  wire [25:0] mem_214_6_W0_addr;
  wire  mem_214_6_W0_clk;
  wire [7:0] mem_214_6_W0_data;
  wire  mem_214_6_W0_en;
  wire  mem_214_6_W0_mask;
  wire [25:0] mem_214_7_R0_addr;
  wire  mem_214_7_R0_clk;
  wire [7:0] mem_214_7_R0_data;
  wire  mem_214_7_R0_en;
  wire [25:0] mem_214_7_W0_addr;
  wire  mem_214_7_W0_clk;
  wire [7:0] mem_214_7_W0_data;
  wire  mem_214_7_W0_en;
  wire  mem_214_7_W0_mask;
  wire [25:0] mem_215_0_R0_addr;
  wire  mem_215_0_R0_clk;
  wire [7:0] mem_215_0_R0_data;
  wire  mem_215_0_R0_en;
  wire [25:0] mem_215_0_W0_addr;
  wire  mem_215_0_W0_clk;
  wire [7:0] mem_215_0_W0_data;
  wire  mem_215_0_W0_en;
  wire  mem_215_0_W0_mask;
  wire [25:0] mem_215_1_R0_addr;
  wire  mem_215_1_R0_clk;
  wire [7:0] mem_215_1_R0_data;
  wire  mem_215_1_R0_en;
  wire [25:0] mem_215_1_W0_addr;
  wire  mem_215_1_W0_clk;
  wire [7:0] mem_215_1_W0_data;
  wire  mem_215_1_W0_en;
  wire  mem_215_1_W0_mask;
  wire [25:0] mem_215_2_R0_addr;
  wire  mem_215_2_R0_clk;
  wire [7:0] mem_215_2_R0_data;
  wire  mem_215_2_R0_en;
  wire [25:0] mem_215_2_W0_addr;
  wire  mem_215_2_W0_clk;
  wire [7:0] mem_215_2_W0_data;
  wire  mem_215_2_W0_en;
  wire  mem_215_2_W0_mask;
  wire [25:0] mem_215_3_R0_addr;
  wire  mem_215_3_R0_clk;
  wire [7:0] mem_215_3_R0_data;
  wire  mem_215_3_R0_en;
  wire [25:0] mem_215_3_W0_addr;
  wire  mem_215_3_W0_clk;
  wire [7:0] mem_215_3_W0_data;
  wire  mem_215_3_W0_en;
  wire  mem_215_3_W0_mask;
  wire [25:0] mem_215_4_R0_addr;
  wire  mem_215_4_R0_clk;
  wire [7:0] mem_215_4_R0_data;
  wire  mem_215_4_R0_en;
  wire [25:0] mem_215_4_W0_addr;
  wire  mem_215_4_W0_clk;
  wire [7:0] mem_215_4_W0_data;
  wire  mem_215_4_W0_en;
  wire  mem_215_4_W0_mask;
  wire [25:0] mem_215_5_R0_addr;
  wire  mem_215_5_R0_clk;
  wire [7:0] mem_215_5_R0_data;
  wire  mem_215_5_R0_en;
  wire [25:0] mem_215_5_W0_addr;
  wire  mem_215_5_W0_clk;
  wire [7:0] mem_215_5_W0_data;
  wire  mem_215_5_W0_en;
  wire  mem_215_5_W0_mask;
  wire [25:0] mem_215_6_R0_addr;
  wire  mem_215_6_R0_clk;
  wire [7:0] mem_215_6_R0_data;
  wire  mem_215_6_R0_en;
  wire [25:0] mem_215_6_W0_addr;
  wire  mem_215_6_W0_clk;
  wire [7:0] mem_215_6_W0_data;
  wire  mem_215_6_W0_en;
  wire  mem_215_6_W0_mask;
  wire [25:0] mem_215_7_R0_addr;
  wire  mem_215_7_R0_clk;
  wire [7:0] mem_215_7_R0_data;
  wire  mem_215_7_R0_en;
  wire [25:0] mem_215_7_W0_addr;
  wire  mem_215_7_W0_clk;
  wire [7:0] mem_215_7_W0_data;
  wire  mem_215_7_W0_en;
  wire  mem_215_7_W0_mask;
  wire [25:0] mem_216_0_R0_addr;
  wire  mem_216_0_R0_clk;
  wire [7:0] mem_216_0_R0_data;
  wire  mem_216_0_R0_en;
  wire [25:0] mem_216_0_W0_addr;
  wire  mem_216_0_W0_clk;
  wire [7:0] mem_216_0_W0_data;
  wire  mem_216_0_W0_en;
  wire  mem_216_0_W0_mask;
  wire [25:0] mem_216_1_R0_addr;
  wire  mem_216_1_R0_clk;
  wire [7:0] mem_216_1_R0_data;
  wire  mem_216_1_R0_en;
  wire [25:0] mem_216_1_W0_addr;
  wire  mem_216_1_W0_clk;
  wire [7:0] mem_216_1_W0_data;
  wire  mem_216_1_W0_en;
  wire  mem_216_1_W0_mask;
  wire [25:0] mem_216_2_R0_addr;
  wire  mem_216_2_R0_clk;
  wire [7:0] mem_216_2_R0_data;
  wire  mem_216_2_R0_en;
  wire [25:0] mem_216_2_W0_addr;
  wire  mem_216_2_W0_clk;
  wire [7:0] mem_216_2_W0_data;
  wire  mem_216_2_W0_en;
  wire  mem_216_2_W0_mask;
  wire [25:0] mem_216_3_R0_addr;
  wire  mem_216_3_R0_clk;
  wire [7:0] mem_216_3_R0_data;
  wire  mem_216_3_R0_en;
  wire [25:0] mem_216_3_W0_addr;
  wire  mem_216_3_W0_clk;
  wire [7:0] mem_216_3_W0_data;
  wire  mem_216_3_W0_en;
  wire  mem_216_3_W0_mask;
  wire [25:0] mem_216_4_R0_addr;
  wire  mem_216_4_R0_clk;
  wire [7:0] mem_216_4_R0_data;
  wire  mem_216_4_R0_en;
  wire [25:0] mem_216_4_W0_addr;
  wire  mem_216_4_W0_clk;
  wire [7:0] mem_216_4_W0_data;
  wire  mem_216_4_W0_en;
  wire  mem_216_4_W0_mask;
  wire [25:0] mem_216_5_R0_addr;
  wire  mem_216_5_R0_clk;
  wire [7:0] mem_216_5_R0_data;
  wire  mem_216_5_R0_en;
  wire [25:0] mem_216_5_W0_addr;
  wire  mem_216_5_W0_clk;
  wire [7:0] mem_216_5_W0_data;
  wire  mem_216_5_W0_en;
  wire  mem_216_5_W0_mask;
  wire [25:0] mem_216_6_R0_addr;
  wire  mem_216_6_R0_clk;
  wire [7:0] mem_216_6_R0_data;
  wire  mem_216_6_R0_en;
  wire [25:0] mem_216_6_W0_addr;
  wire  mem_216_6_W0_clk;
  wire [7:0] mem_216_6_W0_data;
  wire  mem_216_6_W0_en;
  wire  mem_216_6_W0_mask;
  wire [25:0] mem_216_7_R0_addr;
  wire  mem_216_7_R0_clk;
  wire [7:0] mem_216_7_R0_data;
  wire  mem_216_7_R0_en;
  wire [25:0] mem_216_7_W0_addr;
  wire  mem_216_7_W0_clk;
  wire [7:0] mem_216_7_W0_data;
  wire  mem_216_7_W0_en;
  wire  mem_216_7_W0_mask;
  wire [25:0] mem_217_0_R0_addr;
  wire  mem_217_0_R0_clk;
  wire [7:0] mem_217_0_R0_data;
  wire  mem_217_0_R0_en;
  wire [25:0] mem_217_0_W0_addr;
  wire  mem_217_0_W0_clk;
  wire [7:0] mem_217_0_W0_data;
  wire  mem_217_0_W0_en;
  wire  mem_217_0_W0_mask;
  wire [25:0] mem_217_1_R0_addr;
  wire  mem_217_1_R0_clk;
  wire [7:0] mem_217_1_R0_data;
  wire  mem_217_1_R0_en;
  wire [25:0] mem_217_1_W0_addr;
  wire  mem_217_1_W0_clk;
  wire [7:0] mem_217_1_W0_data;
  wire  mem_217_1_W0_en;
  wire  mem_217_1_W0_mask;
  wire [25:0] mem_217_2_R0_addr;
  wire  mem_217_2_R0_clk;
  wire [7:0] mem_217_2_R0_data;
  wire  mem_217_2_R0_en;
  wire [25:0] mem_217_2_W0_addr;
  wire  mem_217_2_W0_clk;
  wire [7:0] mem_217_2_W0_data;
  wire  mem_217_2_W0_en;
  wire  mem_217_2_W0_mask;
  wire [25:0] mem_217_3_R0_addr;
  wire  mem_217_3_R0_clk;
  wire [7:0] mem_217_3_R0_data;
  wire  mem_217_3_R0_en;
  wire [25:0] mem_217_3_W0_addr;
  wire  mem_217_3_W0_clk;
  wire [7:0] mem_217_3_W0_data;
  wire  mem_217_3_W0_en;
  wire  mem_217_3_W0_mask;
  wire [25:0] mem_217_4_R0_addr;
  wire  mem_217_4_R0_clk;
  wire [7:0] mem_217_4_R0_data;
  wire  mem_217_4_R0_en;
  wire [25:0] mem_217_4_W0_addr;
  wire  mem_217_4_W0_clk;
  wire [7:0] mem_217_4_W0_data;
  wire  mem_217_4_W0_en;
  wire  mem_217_4_W0_mask;
  wire [25:0] mem_217_5_R0_addr;
  wire  mem_217_5_R0_clk;
  wire [7:0] mem_217_5_R0_data;
  wire  mem_217_5_R0_en;
  wire [25:0] mem_217_5_W0_addr;
  wire  mem_217_5_W0_clk;
  wire [7:0] mem_217_5_W0_data;
  wire  mem_217_5_W0_en;
  wire  mem_217_5_W0_mask;
  wire [25:0] mem_217_6_R0_addr;
  wire  mem_217_6_R0_clk;
  wire [7:0] mem_217_6_R0_data;
  wire  mem_217_6_R0_en;
  wire [25:0] mem_217_6_W0_addr;
  wire  mem_217_6_W0_clk;
  wire [7:0] mem_217_6_W0_data;
  wire  mem_217_6_W0_en;
  wire  mem_217_6_W0_mask;
  wire [25:0] mem_217_7_R0_addr;
  wire  mem_217_7_R0_clk;
  wire [7:0] mem_217_7_R0_data;
  wire  mem_217_7_R0_en;
  wire [25:0] mem_217_7_W0_addr;
  wire  mem_217_7_W0_clk;
  wire [7:0] mem_217_7_W0_data;
  wire  mem_217_7_W0_en;
  wire  mem_217_7_W0_mask;
  wire [25:0] mem_218_0_R0_addr;
  wire  mem_218_0_R0_clk;
  wire [7:0] mem_218_0_R0_data;
  wire  mem_218_0_R0_en;
  wire [25:0] mem_218_0_W0_addr;
  wire  mem_218_0_W0_clk;
  wire [7:0] mem_218_0_W0_data;
  wire  mem_218_0_W0_en;
  wire  mem_218_0_W0_mask;
  wire [25:0] mem_218_1_R0_addr;
  wire  mem_218_1_R0_clk;
  wire [7:0] mem_218_1_R0_data;
  wire  mem_218_1_R0_en;
  wire [25:0] mem_218_1_W0_addr;
  wire  mem_218_1_W0_clk;
  wire [7:0] mem_218_1_W0_data;
  wire  mem_218_1_W0_en;
  wire  mem_218_1_W0_mask;
  wire [25:0] mem_218_2_R0_addr;
  wire  mem_218_2_R0_clk;
  wire [7:0] mem_218_2_R0_data;
  wire  mem_218_2_R0_en;
  wire [25:0] mem_218_2_W0_addr;
  wire  mem_218_2_W0_clk;
  wire [7:0] mem_218_2_W0_data;
  wire  mem_218_2_W0_en;
  wire  mem_218_2_W0_mask;
  wire [25:0] mem_218_3_R0_addr;
  wire  mem_218_3_R0_clk;
  wire [7:0] mem_218_3_R0_data;
  wire  mem_218_3_R0_en;
  wire [25:0] mem_218_3_W0_addr;
  wire  mem_218_3_W0_clk;
  wire [7:0] mem_218_3_W0_data;
  wire  mem_218_3_W0_en;
  wire  mem_218_3_W0_mask;
  wire [25:0] mem_218_4_R0_addr;
  wire  mem_218_4_R0_clk;
  wire [7:0] mem_218_4_R0_data;
  wire  mem_218_4_R0_en;
  wire [25:0] mem_218_4_W0_addr;
  wire  mem_218_4_W0_clk;
  wire [7:0] mem_218_4_W0_data;
  wire  mem_218_4_W0_en;
  wire  mem_218_4_W0_mask;
  wire [25:0] mem_218_5_R0_addr;
  wire  mem_218_5_R0_clk;
  wire [7:0] mem_218_5_R0_data;
  wire  mem_218_5_R0_en;
  wire [25:0] mem_218_5_W0_addr;
  wire  mem_218_5_W0_clk;
  wire [7:0] mem_218_5_W0_data;
  wire  mem_218_5_W0_en;
  wire  mem_218_5_W0_mask;
  wire [25:0] mem_218_6_R0_addr;
  wire  mem_218_6_R0_clk;
  wire [7:0] mem_218_6_R0_data;
  wire  mem_218_6_R0_en;
  wire [25:0] mem_218_6_W0_addr;
  wire  mem_218_6_W0_clk;
  wire [7:0] mem_218_6_W0_data;
  wire  mem_218_6_W0_en;
  wire  mem_218_6_W0_mask;
  wire [25:0] mem_218_7_R0_addr;
  wire  mem_218_7_R0_clk;
  wire [7:0] mem_218_7_R0_data;
  wire  mem_218_7_R0_en;
  wire [25:0] mem_218_7_W0_addr;
  wire  mem_218_7_W0_clk;
  wire [7:0] mem_218_7_W0_data;
  wire  mem_218_7_W0_en;
  wire  mem_218_7_W0_mask;
  wire [25:0] mem_219_0_R0_addr;
  wire  mem_219_0_R0_clk;
  wire [7:0] mem_219_0_R0_data;
  wire  mem_219_0_R0_en;
  wire [25:0] mem_219_0_W0_addr;
  wire  mem_219_0_W0_clk;
  wire [7:0] mem_219_0_W0_data;
  wire  mem_219_0_W0_en;
  wire  mem_219_0_W0_mask;
  wire [25:0] mem_219_1_R0_addr;
  wire  mem_219_1_R0_clk;
  wire [7:0] mem_219_1_R0_data;
  wire  mem_219_1_R0_en;
  wire [25:0] mem_219_1_W0_addr;
  wire  mem_219_1_W0_clk;
  wire [7:0] mem_219_1_W0_data;
  wire  mem_219_1_W0_en;
  wire  mem_219_1_W0_mask;
  wire [25:0] mem_219_2_R0_addr;
  wire  mem_219_2_R0_clk;
  wire [7:0] mem_219_2_R0_data;
  wire  mem_219_2_R0_en;
  wire [25:0] mem_219_2_W0_addr;
  wire  mem_219_2_W0_clk;
  wire [7:0] mem_219_2_W0_data;
  wire  mem_219_2_W0_en;
  wire  mem_219_2_W0_mask;
  wire [25:0] mem_219_3_R0_addr;
  wire  mem_219_3_R0_clk;
  wire [7:0] mem_219_3_R0_data;
  wire  mem_219_3_R0_en;
  wire [25:0] mem_219_3_W0_addr;
  wire  mem_219_3_W0_clk;
  wire [7:0] mem_219_3_W0_data;
  wire  mem_219_3_W0_en;
  wire  mem_219_3_W0_mask;
  wire [25:0] mem_219_4_R0_addr;
  wire  mem_219_4_R0_clk;
  wire [7:0] mem_219_4_R0_data;
  wire  mem_219_4_R0_en;
  wire [25:0] mem_219_4_W0_addr;
  wire  mem_219_4_W0_clk;
  wire [7:0] mem_219_4_W0_data;
  wire  mem_219_4_W0_en;
  wire  mem_219_4_W0_mask;
  wire [25:0] mem_219_5_R0_addr;
  wire  mem_219_5_R0_clk;
  wire [7:0] mem_219_5_R0_data;
  wire  mem_219_5_R0_en;
  wire [25:0] mem_219_5_W0_addr;
  wire  mem_219_5_W0_clk;
  wire [7:0] mem_219_5_W0_data;
  wire  mem_219_5_W0_en;
  wire  mem_219_5_W0_mask;
  wire [25:0] mem_219_6_R0_addr;
  wire  mem_219_6_R0_clk;
  wire [7:0] mem_219_6_R0_data;
  wire  mem_219_6_R0_en;
  wire [25:0] mem_219_6_W0_addr;
  wire  mem_219_6_W0_clk;
  wire [7:0] mem_219_6_W0_data;
  wire  mem_219_6_W0_en;
  wire  mem_219_6_W0_mask;
  wire [25:0] mem_219_7_R0_addr;
  wire  mem_219_7_R0_clk;
  wire [7:0] mem_219_7_R0_data;
  wire  mem_219_7_R0_en;
  wire [25:0] mem_219_7_W0_addr;
  wire  mem_219_7_W0_clk;
  wire [7:0] mem_219_7_W0_data;
  wire  mem_219_7_W0_en;
  wire  mem_219_7_W0_mask;
  wire [25:0] mem_220_0_R0_addr;
  wire  mem_220_0_R0_clk;
  wire [7:0] mem_220_0_R0_data;
  wire  mem_220_0_R0_en;
  wire [25:0] mem_220_0_W0_addr;
  wire  mem_220_0_W0_clk;
  wire [7:0] mem_220_0_W0_data;
  wire  mem_220_0_W0_en;
  wire  mem_220_0_W0_mask;
  wire [25:0] mem_220_1_R0_addr;
  wire  mem_220_1_R0_clk;
  wire [7:0] mem_220_1_R0_data;
  wire  mem_220_1_R0_en;
  wire [25:0] mem_220_1_W0_addr;
  wire  mem_220_1_W0_clk;
  wire [7:0] mem_220_1_W0_data;
  wire  mem_220_1_W0_en;
  wire  mem_220_1_W0_mask;
  wire [25:0] mem_220_2_R0_addr;
  wire  mem_220_2_R0_clk;
  wire [7:0] mem_220_2_R0_data;
  wire  mem_220_2_R0_en;
  wire [25:0] mem_220_2_W0_addr;
  wire  mem_220_2_W0_clk;
  wire [7:0] mem_220_2_W0_data;
  wire  mem_220_2_W0_en;
  wire  mem_220_2_W0_mask;
  wire [25:0] mem_220_3_R0_addr;
  wire  mem_220_3_R0_clk;
  wire [7:0] mem_220_3_R0_data;
  wire  mem_220_3_R0_en;
  wire [25:0] mem_220_3_W0_addr;
  wire  mem_220_3_W0_clk;
  wire [7:0] mem_220_3_W0_data;
  wire  mem_220_3_W0_en;
  wire  mem_220_3_W0_mask;
  wire [25:0] mem_220_4_R0_addr;
  wire  mem_220_4_R0_clk;
  wire [7:0] mem_220_4_R0_data;
  wire  mem_220_4_R0_en;
  wire [25:0] mem_220_4_W0_addr;
  wire  mem_220_4_W0_clk;
  wire [7:0] mem_220_4_W0_data;
  wire  mem_220_4_W0_en;
  wire  mem_220_4_W0_mask;
  wire [25:0] mem_220_5_R0_addr;
  wire  mem_220_5_R0_clk;
  wire [7:0] mem_220_5_R0_data;
  wire  mem_220_5_R0_en;
  wire [25:0] mem_220_5_W0_addr;
  wire  mem_220_5_W0_clk;
  wire [7:0] mem_220_5_W0_data;
  wire  mem_220_5_W0_en;
  wire  mem_220_5_W0_mask;
  wire [25:0] mem_220_6_R0_addr;
  wire  mem_220_6_R0_clk;
  wire [7:0] mem_220_6_R0_data;
  wire  mem_220_6_R0_en;
  wire [25:0] mem_220_6_W0_addr;
  wire  mem_220_6_W0_clk;
  wire [7:0] mem_220_6_W0_data;
  wire  mem_220_6_W0_en;
  wire  mem_220_6_W0_mask;
  wire [25:0] mem_220_7_R0_addr;
  wire  mem_220_7_R0_clk;
  wire [7:0] mem_220_7_R0_data;
  wire  mem_220_7_R0_en;
  wire [25:0] mem_220_7_W0_addr;
  wire  mem_220_7_W0_clk;
  wire [7:0] mem_220_7_W0_data;
  wire  mem_220_7_W0_en;
  wire  mem_220_7_W0_mask;
  wire [25:0] mem_221_0_R0_addr;
  wire  mem_221_0_R0_clk;
  wire [7:0] mem_221_0_R0_data;
  wire  mem_221_0_R0_en;
  wire [25:0] mem_221_0_W0_addr;
  wire  mem_221_0_W0_clk;
  wire [7:0] mem_221_0_W0_data;
  wire  mem_221_0_W0_en;
  wire  mem_221_0_W0_mask;
  wire [25:0] mem_221_1_R0_addr;
  wire  mem_221_1_R0_clk;
  wire [7:0] mem_221_1_R0_data;
  wire  mem_221_1_R0_en;
  wire [25:0] mem_221_1_W0_addr;
  wire  mem_221_1_W0_clk;
  wire [7:0] mem_221_1_W0_data;
  wire  mem_221_1_W0_en;
  wire  mem_221_1_W0_mask;
  wire [25:0] mem_221_2_R0_addr;
  wire  mem_221_2_R0_clk;
  wire [7:0] mem_221_2_R0_data;
  wire  mem_221_2_R0_en;
  wire [25:0] mem_221_2_W0_addr;
  wire  mem_221_2_W0_clk;
  wire [7:0] mem_221_2_W0_data;
  wire  mem_221_2_W0_en;
  wire  mem_221_2_W0_mask;
  wire [25:0] mem_221_3_R0_addr;
  wire  mem_221_3_R0_clk;
  wire [7:0] mem_221_3_R0_data;
  wire  mem_221_3_R0_en;
  wire [25:0] mem_221_3_W0_addr;
  wire  mem_221_3_W0_clk;
  wire [7:0] mem_221_3_W0_data;
  wire  mem_221_3_W0_en;
  wire  mem_221_3_W0_mask;
  wire [25:0] mem_221_4_R0_addr;
  wire  mem_221_4_R0_clk;
  wire [7:0] mem_221_4_R0_data;
  wire  mem_221_4_R0_en;
  wire [25:0] mem_221_4_W0_addr;
  wire  mem_221_4_W0_clk;
  wire [7:0] mem_221_4_W0_data;
  wire  mem_221_4_W0_en;
  wire  mem_221_4_W0_mask;
  wire [25:0] mem_221_5_R0_addr;
  wire  mem_221_5_R0_clk;
  wire [7:0] mem_221_5_R0_data;
  wire  mem_221_5_R0_en;
  wire [25:0] mem_221_5_W0_addr;
  wire  mem_221_5_W0_clk;
  wire [7:0] mem_221_5_W0_data;
  wire  mem_221_5_W0_en;
  wire  mem_221_5_W0_mask;
  wire [25:0] mem_221_6_R0_addr;
  wire  mem_221_6_R0_clk;
  wire [7:0] mem_221_6_R0_data;
  wire  mem_221_6_R0_en;
  wire [25:0] mem_221_6_W0_addr;
  wire  mem_221_6_W0_clk;
  wire [7:0] mem_221_6_W0_data;
  wire  mem_221_6_W0_en;
  wire  mem_221_6_W0_mask;
  wire [25:0] mem_221_7_R0_addr;
  wire  mem_221_7_R0_clk;
  wire [7:0] mem_221_7_R0_data;
  wire  mem_221_7_R0_en;
  wire [25:0] mem_221_7_W0_addr;
  wire  mem_221_7_W0_clk;
  wire [7:0] mem_221_7_W0_data;
  wire  mem_221_7_W0_en;
  wire  mem_221_7_W0_mask;
  wire [25:0] mem_222_0_R0_addr;
  wire  mem_222_0_R0_clk;
  wire [7:0] mem_222_0_R0_data;
  wire  mem_222_0_R0_en;
  wire [25:0] mem_222_0_W0_addr;
  wire  mem_222_0_W0_clk;
  wire [7:0] mem_222_0_W0_data;
  wire  mem_222_0_W0_en;
  wire  mem_222_0_W0_mask;
  wire [25:0] mem_222_1_R0_addr;
  wire  mem_222_1_R0_clk;
  wire [7:0] mem_222_1_R0_data;
  wire  mem_222_1_R0_en;
  wire [25:0] mem_222_1_W0_addr;
  wire  mem_222_1_W0_clk;
  wire [7:0] mem_222_1_W0_data;
  wire  mem_222_1_W0_en;
  wire  mem_222_1_W0_mask;
  wire [25:0] mem_222_2_R0_addr;
  wire  mem_222_2_R0_clk;
  wire [7:0] mem_222_2_R0_data;
  wire  mem_222_2_R0_en;
  wire [25:0] mem_222_2_W0_addr;
  wire  mem_222_2_W0_clk;
  wire [7:0] mem_222_2_W0_data;
  wire  mem_222_2_W0_en;
  wire  mem_222_2_W0_mask;
  wire [25:0] mem_222_3_R0_addr;
  wire  mem_222_3_R0_clk;
  wire [7:0] mem_222_3_R0_data;
  wire  mem_222_3_R0_en;
  wire [25:0] mem_222_3_W0_addr;
  wire  mem_222_3_W0_clk;
  wire [7:0] mem_222_3_W0_data;
  wire  mem_222_3_W0_en;
  wire  mem_222_3_W0_mask;
  wire [25:0] mem_222_4_R0_addr;
  wire  mem_222_4_R0_clk;
  wire [7:0] mem_222_4_R0_data;
  wire  mem_222_4_R0_en;
  wire [25:0] mem_222_4_W0_addr;
  wire  mem_222_4_W0_clk;
  wire [7:0] mem_222_4_W0_data;
  wire  mem_222_4_W0_en;
  wire  mem_222_4_W0_mask;
  wire [25:0] mem_222_5_R0_addr;
  wire  mem_222_5_R0_clk;
  wire [7:0] mem_222_5_R0_data;
  wire  mem_222_5_R0_en;
  wire [25:0] mem_222_5_W0_addr;
  wire  mem_222_5_W0_clk;
  wire [7:0] mem_222_5_W0_data;
  wire  mem_222_5_W0_en;
  wire  mem_222_5_W0_mask;
  wire [25:0] mem_222_6_R0_addr;
  wire  mem_222_6_R0_clk;
  wire [7:0] mem_222_6_R0_data;
  wire  mem_222_6_R0_en;
  wire [25:0] mem_222_6_W0_addr;
  wire  mem_222_6_W0_clk;
  wire [7:0] mem_222_6_W0_data;
  wire  mem_222_6_W0_en;
  wire  mem_222_6_W0_mask;
  wire [25:0] mem_222_7_R0_addr;
  wire  mem_222_7_R0_clk;
  wire [7:0] mem_222_7_R0_data;
  wire  mem_222_7_R0_en;
  wire [25:0] mem_222_7_W0_addr;
  wire  mem_222_7_W0_clk;
  wire [7:0] mem_222_7_W0_data;
  wire  mem_222_7_W0_en;
  wire  mem_222_7_W0_mask;
  wire [25:0] mem_223_0_R0_addr;
  wire  mem_223_0_R0_clk;
  wire [7:0] mem_223_0_R0_data;
  wire  mem_223_0_R0_en;
  wire [25:0] mem_223_0_W0_addr;
  wire  mem_223_0_W0_clk;
  wire [7:0] mem_223_0_W0_data;
  wire  mem_223_0_W0_en;
  wire  mem_223_0_W0_mask;
  wire [25:0] mem_223_1_R0_addr;
  wire  mem_223_1_R0_clk;
  wire [7:0] mem_223_1_R0_data;
  wire  mem_223_1_R0_en;
  wire [25:0] mem_223_1_W0_addr;
  wire  mem_223_1_W0_clk;
  wire [7:0] mem_223_1_W0_data;
  wire  mem_223_1_W0_en;
  wire  mem_223_1_W0_mask;
  wire [25:0] mem_223_2_R0_addr;
  wire  mem_223_2_R0_clk;
  wire [7:0] mem_223_2_R0_data;
  wire  mem_223_2_R0_en;
  wire [25:0] mem_223_2_W0_addr;
  wire  mem_223_2_W0_clk;
  wire [7:0] mem_223_2_W0_data;
  wire  mem_223_2_W0_en;
  wire  mem_223_2_W0_mask;
  wire [25:0] mem_223_3_R0_addr;
  wire  mem_223_3_R0_clk;
  wire [7:0] mem_223_3_R0_data;
  wire  mem_223_3_R0_en;
  wire [25:0] mem_223_3_W0_addr;
  wire  mem_223_3_W0_clk;
  wire [7:0] mem_223_3_W0_data;
  wire  mem_223_3_W0_en;
  wire  mem_223_3_W0_mask;
  wire [25:0] mem_223_4_R0_addr;
  wire  mem_223_4_R0_clk;
  wire [7:0] mem_223_4_R0_data;
  wire  mem_223_4_R0_en;
  wire [25:0] mem_223_4_W0_addr;
  wire  mem_223_4_W0_clk;
  wire [7:0] mem_223_4_W0_data;
  wire  mem_223_4_W0_en;
  wire  mem_223_4_W0_mask;
  wire [25:0] mem_223_5_R0_addr;
  wire  mem_223_5_R0_clk;
  wire [7:0] mem_223_5_R0_data;
  wire  mem_223_5_R0_en;
  wire [25:0] mem_223_5_W0_addr;
  wire  mem_223_5_W0_clk;
  wire [7:0] mem_223_5_W0_data;
  wire  mem_223_5_W0_en;
  wire  mem_223_5_W0_mask;
  wire [25:0] mem_223_6_R0_addr;
  wire  mem_223_6_R0_clk;
  wire [7:0] mem_223_6_R0_data;
  wire  mem_223_6_R0_en;
  wire [25:0] mem_223_6_W0_addr;
  wire  mem_223_6_W0_clk;
  wire [7:0] mem_223_6_W0_data;
  wire  mem_223_6_W0_en;
  wire  mem_223_6_W0_mask;
  wire [25:0] mem_223_7_R0_addr;
  wire  mem_223_7_R0_clk;
  wire [7:0] mem_223_7_R0_data;
  wire  mem_223_7_R0_en;
  wire [25:0] mem_223_7_W0_addr;
  wire  mem_223_7_W0_clk;
  wire [7:0] mem_223_7_W0_data;
  wire  mem_223_7_W0_en;
  wire  mem_223_7_W0_mask;
  wire [25:0] mem_224_0_R0_addr;
  wire  mem_224_0_R0_clk;
  wire [7:0] mem_224_0_R0_data;
  wire  mem_224_0_R0_en;
  wire [25:0] mem_224_0_W0_addr;
  wire  mem_224_0_W0_clk;
  wire [7:0] mem_224_0_W0_data;
  wire  mem_224_0_W0_en;
  wire  mem_224_0_W0_mask;
  wire [25:0] mem_224_1_R0_addr;
  wire  mem_224_1_R0_clk;
  wire [7:0] mem_224_1_R0_data;
  wire  mem_224_1_R0_en;
  wire [25:0] mem_224_1_W0_addr;
  wire  mem_224_1_W0_clk;
  wire [7:0] mem_224_1_W0_data;
  wire  mem_224_1_W0_en;
  wire  mem_224_1_W0_mask;
  wire [25:0] mem_224_2_R0_addr;
  wire  mem_224_2_R0_clk;
  wire [7:0] mem_224_2_R0_data;
  wire  mem_224_2_R0_en;
  wire [25:0] mem_224_2_W0_addr;
  wire  mem_224_2_W0_clk;
  wire [7:0] mem_224_2_W0_data;
  wire  mem_224_2_W0_en;
  wire  mem_224_2_W0_mask;
  wire [25:0] mem_224_3_R0_addr;
  wire  mem_224_3_R0_clk;
  wire [7:0] mem_224_3_R0_data;
  wire  mem_224_3_R0_en;
  wire [25:0] mem_224_3_W0_addr;
  wire  mem_224_3_W0_clk;
  wire [7:0] mem_224_3_W0_data;
  wire  mem_224_3_W0_en;
  wire  mem_224_3_W0_mask;
  wire [25:0] mem_224_4_R0_addr;
  wire  mem_224_4_R0_clk;
  wire [7:0] mem_224_4_R0_data;
  wire  mem_224_4_R0_en;
  wire [25:0] mem_224_4_W0_addr;
  wire  mem_224_4_W0_clk;
  wire [7:0] mem_224_4_W0_data;
  wire  mem_224_4_W0_en;
  wire  mem_224_4_W0_mask;
  wire [25:0] mem_224_5_R0_addr;
  wire  mem_224_5_R0_clk;
  wire [7:0] mem_224_5_R0_data;
  wire  mem_224_5_R0_en;
  wire [25:0] mem_224_5_W0_addr;
  wire  mem_224_5_W0_clk;
  wire [7:0] mem_224_5_W0_data;
  wire  mem_224_5_W0_en;
  wire  mem_224_5_W0_mask;
  wire [25:0] mem_224_6_R0_addr;
  wire  mem_224_6_R0_clk;
  wire [7:0] mem_224_6_R0_data;
  wire  mem_224_6_R0_en;
  wire [25:0] mem_224_6_W0_addr;
  wire  mem_224_6_W0_clk;
  wire [7:0] mem_224_6_W0_data;
  wire  mem_224_6_W0_en;
  wire  mem_224_6_W0_mask;
  wire [25:0] mem_224_7_R0_addr;
  wire  mem_224_7_R0_clk;
  wire [7:0] mem_224_7_R0_data;
  wire  mem_224_7_R0_en;
  wire [25:0] mem_224_7_W0_addr;
  wire  mem_224_7_W0_clk;
  wire [7:0] mem_224_7_W0_data;
  wire  mem_224_7_W0_en;
  wire  mem_224_7_W0_mask;
  wire [25:0] mem_225_0_R0_addr;
  wire  mem_225_0_R0_clk;
  wire [7:0] mem_225_0_R0_data;
  wire  mem_225_0_R0_en;
  wire [25:0] mem_225_0_W0_addr;
  wire  mem_225_0_W0_clk;
  wire [7:0] mem_225_0_W0_data;
  wire  mem_225_0_W0_en;
  wire  mem_225_0_W0_mask;
  wire [25:0] mem_225_1_R0_addr;
  wire  mem_225_1_R0_clk;
  wire [7:0] mem_225_1_R0_data;
  wire  mem_225_1_R0_en;
  wire [25:0] mem_225_1_W0_addr;
  wire  mem_225_1_W0_clk;
  wire [7:0] mem_225_1_W0_data;
  wire  mem_225_1_W0_en;
  wire  mem_225_1_W0_mask;
  wire [25:0] mem_225_2_R0_addr;
  wire  mem_225_2_R0_clk;
  wire [7:0] mem_225_2_R0_data;
  wire  mem_225_2_R0_en;
  wire [25:0] mem_225_2_W0_addr;
  wire  mem_225_2_W0_clk;
  wire [7:0] mem_225_2_W0_data;
  wire  mem_225_2_W0_en;
  wire  mem_225_2_W0_mask;
  wire [25:0] mem_225_3_R0_addr;
  wire  mem_225_3_R0_clk;
  wire [7:0] mem_225_3_R0_data;
  wire  mem_225_3_R0_en;
  wire [25:0] mem_225_3_W0_addr;
  wire  mem_225_3_W0_clk;
  wire [7:0] mem_225_3_W0_data;
  wire  mem_225_3_W0_en;
  wire  mem_225_3_W0_mask;
  wire [25:0] mem_225_4_R0_addr;
  wire  mem_225_4_R0_clk;
  wire [7:0] mem_225_4_R0_data;
  wire  mem_225_4_R0_en;
  wire [25:0] mem_225_4_W0_addr;
  wire  mem_225_4_W0_clk;
  wire [7:0] mem_225_4_W0_data;
  wire  mem_225_4_W0_en;
  wire  mem_225_4_W0_mask;
  wire [25:0] mem_225_5_R0_addr;
  wire  mem_225_5_R0_clk;
  wire [7:0] mem_225_5_R0_data;
  wire  mem_225_5_R0_en;
  wire [25:0] mem_225_5_W0_addr;
  wire  mem_225_5_W0_clk;
  wire [7:0] mem_225_5_W0_data;
  wire  mem_225_5_W0_en;
  wire  mem_225_5_W0_mask;
  wire [25:0] mem_225_6_R0_addr;
  wire  mem_225_6_R0_clk;
  wire [7:0] mem_225_6_R0_data;
  wire  mem_225_6_R0_en;
  wire [25:0] mem_225_6_W0_addr;
  wire  mem_225_6_W0_clk;
  wire [7:0] mem_225_6_W0_data;
  wire  mem_225_6_W0_en;
  wire  mem_225_6_W0_mask;
  wire [25:0] mem_225_7_R0_addr;
  wire  mem_225_7_R0_clk;
  wire [7:0] mem_225_7_R0_data;
  wire  mem_225_7_R0_en;
  wire [25:0] mem_225_7_W0_addr;
  wire  mem_225_7_W0_clk;
  wire [7:0] mem_225_7_W0_data;
  wire  mem_225_7_W0_en;
  wire  mem_225_7_W0_mask;
  wire [25:0] mem_226_0_R0_addr;
  wire  mem_226_0_R0_clk;
  wire [7:0] mem_226_0_R0_data;
  wire  mem_226_0_R0_en;
  wire [25:0] mem_226_0_W0_addr;
  wire  mem_226_0_W0_clk;
  wire [7:0] mem_226_0_W0_data;
  wire  mem_226_0_W0_en;
  wire  mem_226_0_W0_mask;
  wire [25:0] mem_226_1_R0_addr;
  wire  mem_226_1_R0_clk;
  wire [7:0] mem_226_1_R0_data;
  wire  mem_226_1_R0_en;
  wire [25:0] mem_226_1_W0_addr;
  wire  mem_226_1_W0_clk;
  wire [7:0] mem_226_1_W0_data;
  wire  mem_226_1_W0_en;
  wire  mem_226_1_W0_mask;
  wire [25:0] mem_226_2_R0_addr;
  wire  mem_226_2_R0_clk;
  wire [7:0] mem_226_2_R0_data;
  wire  mem_226_2_R0_en;
  wire [25:0] mem_226_2_W0_addr;
  wire  mem_226_2_W0_clk;
  wire [7:0] mem_226_2_W0_data;
  wire  mem_226_2_W0_en;
  wire  mem_226_2_W0_mask;
  wire [25:0] mem_226_3_R0_addr;
  wire  mem_226_3_R0_clk;
  wire [7:0] mem_226_3_R0_data;
  wire  mem_226_3_R0_en;
  wire [25:0] mem_226_3_W0_addr;
  wire  mem_226_3_W0_clk;
  wire [7:0] mem_226_3_W0_data;
  wire  mem_226_3_W0_en;
  wire  mem_226_3_W0_mask;
  wire [25:0] mem_226_4_R0_addr;
  wire  mem_226_4_R0_clk;
  wire [7:0] mem_226_4_R0_data;
  wire  mem_226_4_R0_en;
  wire [25:0] mem_226_4_W0_addr;
  wire  mem_226_4_W0_clk;
  wire [7:0] mem_226_4_W0_data;
  wire  mem_226_4_W0_en;
  wire  mem_226_4_W0_mask;
  wire [25:0] mem_226_5_R0_addr;
  wire  mem_226_5_R0_clk;
  wire [7:0] mem_226_5_R0_data;
  wire  mem_226_5_R0_en;
  wire [25:0] mem_226_5_W0_addr;
  wire  mem_226_5_W0_clk;
  wire [7:0] mem_226_5_W0_data;
  wire  mem_226_5_W0_en;
  wire  mem_226_5_W0_mask;
  wire [25:0] mem_226_6_R0_addr;
  wire  mem_226_6_R0_clk;
  wire [7:0] mem_226_6_R0_data;
  wire  mem_226_6_R0_en;
  wire [25:0] mem_226_6_W0_addr;
  wire  mem_226_6_W0_clk;
  wire [7:0] mem_226_6_W0_data;
  wire  mem_226_6_W0_en;
  wire  mem_226_6_W0_mask;
  wire [25:0] mem_226_7_R0_addr;
  wire  mem_226_7_R0_clk;
  wire [7:0] mem_226_7_R0_data;
  wire  mem_226_7_R0_en;
  wire [25:0] mem_226_7_W0_addr;
  wire  mem_226_7_W0_clk;
  wire [7:0] mem_226_7_W0_data;
  wire  mem_226_7_W0_en;
  wire  mem_226_7_W0_mask;
  wire [25:0] mem_227_0_R0_addr;
  wire  mem_227_0_R0_clk;
  wire [7:0] mem_227_0_R0_data;
  wire  mem_227_0_R0_en;
  wire [25:0] mem_227_0_W0_addr;
  wire  mem_227_0_W0_clk;
  wire [7:0] mem_227_0_W0_data;
  wire  mem_227_0_W0_en;
  wire  mem_227_0_W0_mask;
  wire [25:0] mem_227_1_R0_addr;
  wire  mem_227_1_R0_clk;
  wire [7:0] mem_227_1_R0_data;
  wire  mem_227_1_R0_en;
  wire [25:0] mem_227_1_W0_addr;
  wire  mem_227_1_W0_clk;
  wire [7:0] mem_227_1_W0_data;
  wire  mem_227_1_W0_en;
  wire  mem_227_1_W0_mask;
  wire [25:0] mem_227_2_R0_addr;
  wire  mem_227_2_R0_clk;
  wire [7:0] mem_227_2_R0_data;
  wire  mem_227_2_R0_en;
  wire [25:0] mem_227_2_W0_addr;
  wire  mem_227_2_W0_clk;
  wire [7:0] mem_227_2_W0_data;
  wire  mem_227_2_W0_en;
  wire  mem_227_2_W0_mask;
  wire [25:0] mem_227_3_R0_addr;
  wire  mem_227_3_R0_clk;
  wire [7:0] mem_227_3_R0_data;
  wire  mem_227_3_R0_en;
  wire [25:0] mem_227_3_W0_addr;
  wire  mem_227_3_W0_clk;
  wire [7:0] mem_227_3_W0_data;
  wire  mem_227_3_W0_en;
  wire  mem_227_3_W0_mask;
  wire [25:0] mem_227_4_R0_addr;
  wire  mem_227_4_R0_clk;
  wire [7:0] mem_227_4_R0_data;
  wire  mem_227_4_R0_en;
  wire [25:0] mem_227_4_W0_addr;
  wire  mem_227_4_W0_clk;
  wire [7:0] mem_227_4_W0_data;
  wire  mem_227_4_W0_en;
  wire  mem_227_4_W0_mask;
  wire [25:0] mem_227_5_R0_addr;
  wire  mem_227_5_R0_clk;
  wire [7:0] mem_227_5_R0_data;
  wire  mem_227_5_R0_en;
  wire [25:0] mem_227_5_W0_addr;
  wire  mem_227_5_W0_clk;
  wire [7:0] mem_227_5_W0_data;
  wire  mem_227_5_W0_en;
  wire  mem_227_5_W0_mask;
  wire [25:0] mem_227_6_R0_addr;
  wire  mem_227_6_R0_clk;
  wire [7:0] mem_227_6_R0_data;
  wire  mem_227_6_R0_en;
  wire [25:0] mem_227_6_W0_addr;
  wire  mem_227_6_W0_clk;
  wire [7:0] mem_227_6_W0_data;
  wire  mem_227_6_W0_en;
  wire  mem_227_6_W0_mask;
  wire [25:0] mem_227_7_R0_addr;
  wire  mem_227_7_R0_clk;
  wire [7:0] mem_227_7_R0_data;
  wire  mem_227_7_R0_en;
  wire [25:0] mem_227_7_W0_addr;
  wire  mem_227_7_W0_clk;
  wire [7:0] mem_227_7_W0_data;
  wire  mem_227_7_W0_en;
  wire  mem_227_7_W0_mask;
  wire [25:0] mem_228_0_R0_addr;
  wire  mem_228_0_R0_clk;
  wire [7:0] mem_228_0_R0_data;
  wire  mem_228_0_R0_en;
  wire [25:0] mem_228_0_W0_addr;
  wire  mem_228_0_W0_clk;
  wire [7:0] mem_228_0_W0_data;
  wire  mem_228_0_W0_en;
  wire  mem_228_0_W0_mask;
  wire [25:0] mem_228_1_R0_addr;
  wire  mem_228_1_R0_clk;
  wire [7:0] mem_228_1_R0_data;
  wire  mem_228_1_R0_en;
  wire [25:0] mem_228_1_W0_addr;
  wire  mem_228_1_W0_clk;
  wire [7:0] mem_228_1_W0_data;
  wire  mem_228_1_W0_en;
  wire  mem_228_1_W0_mask;
  wire [25:0] mem_228_2_R0_addr;
  wire  mem_228_2_R0_clk;
  wire [7:0] mem_228_2_R0_data;
  wire  mem_228_2_R0_en;
  wire [25:0] mem_228_2_W0_addr;
  wire  mem_228_2_W0_clk;
  wire [7:0] mem_228_2_W0_data;
  wire  mem_228_2_W0_en;
  wire  mem_228_2_W0_mask;
  wire [25:0] mem_228_3_R0_addr;
  wire  mem_228_3_R0_clk;
  wire [7:0] mem_228_3_R0_data;
  wire  mem_228_3_R0_en;
  wire [25:0] mem_228_3_W0_addr;
  wire  mem_228_3_W0_clk;
  wire [7:0] mem_228_3_W0_data;
  wire  mem_228_3_W0_en;
  wire  mem_228_3_W0_mask;
  wire [25:0] mem_228_4_R0_addr;
  wire  mem_228_4_R0_clk;
  wire [7:0] mem_228_4_R0_data;
  wire  mem_228_4_R0_en;
  wire [25:0] mem_228_4_W0_addr;
  wire  mem_228_4_W0_clk;
  wire [7:0] mem_228_4_W0_data;
  wire  mem_228_4_W0_en;
  wire  mem_228_4_W0_mask;
  wire [25:0] mem_228_5_R0_addr;
  wire  mem_228_5_R0_clk;
  wire [7:0] mem_228_5_R0_data;
  wire  mem_228_5_R0_en;
  wire [25:0] mem_228_5_W0_addr;
  wire  mem_228_5_W0_clk;
  wire [7:0] mem_228_5_W0_data;
  wire  mem_228_5_W0_en;
  wire  mem_228_5_W0_mask;
  wire [25:0] mem_228_6_R0_addr;
  wire  mem_228_6_R0_clk;
  wire [7:0] mem_228_6_R0_data;
  wire  mem_228_6_R0_en;
  wire [25:0] mem_228_6_W0_addr;
  wire  mem_228_6_W0_clk;
  wire [7:0] mem_228_6_W0_data;
  wire  mem_228_6_W0_en;
  wire  mem_228_6_W0_mask;
  wire [25:0] mem_228_7_R0_addr;
  wire  mem_228_7_R0_clk;
  wire [7:0] mem_228_7_R0_data;
  wire  mem_228_7_R0_en;
  wire [25:0] mem_228_7_W0_addr;
  wire  mem_228_7_W0_clk;
  wire [7:0] mem_228_7_W0_data;
  wire  mem_228_7_W0_en;
  wire  mem_228_7_W0_mask;
  wire [25:0] mem_229_0_R0_addr;
  wire  mem_229_0_R0_clk;
  wire [7:0] mem_229_0_R0_data;
  wire  mem_229_0_R0_en;
  wire [25:0] mem_229_0_W0_addr;
  wire  mem_229_0_W0_clk;
  wire [7:0] mem_229_0_W0_data;
  wire  mem_229_0_W0_en;
  wire  mem_229_0_W0_mask;
  wire [25:0] mem_229_1_R0_addr;
  wire  mem_229_1_R0_clk;
  wire [7:0] mem_229_1_R0_data;
  wire  mem_229_1_R0_en;
  wire [25:0] mem_229_1_W0_addr;
  wire  mem_229_1_W0_clk;
  wire [7:0] mem_229_1_W0_data;
  wire  mem_229_1_W0_en;
  wire  mem_229_1_W0_mask;
  wire [25:0] mem_229_2_R0_addr;
  wire  mem_229_2_R0_clk;
  wire [7:0] mem_229_2_R0_data;
  wire  mem_229_2_R0_en;
  wire [25:0] mem_229_2_W0_addr;
  wire  mem_229_2_W0_clk;
  wire [7:0] mem_229_2_W0_data;
  wire  mem_229_2_W0_en;
  wire  mem_229_2_W0_mask;
  wire [25:0] mem_229_3_R0_addr;
  wire  mem_229_3_R0_clk;
  wire [7:0] mem_229_3_R0_data;
  wire  mem_229_3_R0_en;
  wire [25:0] mem_229_3_W0_addr;
  wire  mem_229_3_W0_clk;
  wire [7:0] mem_229_3_W0_data;
  wire  mem_229_3_W0_en;
  wire  mem_229_3_W0_mask;
  wire [25:0] mem_229_4_R0_addr;
  wire  mem_229_4_R0_clk;
  wire [7:0] mem_229_4_R0_data;
  wire  mem_229_4_R0_en;
  wire [25:0] mem_229_4_W0_addr;
  wire  mem_229_4_W0_clk;
  wire [7:0] mem_229_4_W0_data;
  wire  mem_229_4_W0_en;
  wire  mem_229_4_W0_mask;
  wire [25:0] mem_229_5_R0_addr;
  wire  mem_229_5_R0_clk;
  wire [7:0] mem_229_5_R0_data;
  wire  mem_229_5_R0_en;
  wire [25:0] mem_229_5_W0_addr;
  wire  mem_229_5_W0_clk;
  wire [7:0] mem_229_5_W0_data;
  wire  mem_229_5_W0_en;
  wire  mem_229_5_W0_mask;
  wire [25:0] mem_229_6_R0_addr;
  wire  mem_229_6_R0_clk;
  wire [7:0] mem_229_6_R0_data;
  wire  mem_229_6_R0_en;
  wire [25:0] mem_229_6_W0_addr;
  wire  mem_229_6_W0_clk;
  wire [7:0] mem_229_6_W0_data;
  wire  mem_229_6_W0_en;
  wire  mem_229_6_W0_mask;
  wire [25:0] mem_229_7_R0_addr;
  wire  mem_229_7_R0_clk;
  wire [7:0] mem_229_7_R0_data;
  wire  mem_229_7_R0_en;
  wire [25:0] mem_229_7_W0_addr;
  wire  mem_229_7_W0_clk;
  wire [7:0] mem_229_7_W0_data;
  wire  mem_229_7_W0_en;
  wire  mem_229_7_W0_mask;
  wire [25:0] mem_230_0_R0_addr;
  wire  mem_230_0_R0_clk;
  wire [7:0] mem_230_0_R0_data;
  wire  mem_230_0_R0_en;
  wire [25:0] mem_230_0_W0_addr;
  wire  mem_230_0_W0_clk;
  wire [7:0] mem_230_0_W0_data;
  wire  mem_230_0_W0_en;
  wire  mem_230_0_W0_mask;
  wire [25:0] mem_230_1_R0_addr;
  wire  mem_230_1_R0_clk;
  wire [7:0] mem_230_1_R0_data;
  wire  mem_230_1_R0_en;
  wire [25:0] mem_230_1_W0_addr;
  wire  mem_230_1_W0_clk;
  wire [7:0] mem_230_1_W0_data;
  wire  mem_230_1_W0_en;
  wire  mem_230_1_W0_mask;
  wire [25:0] mem_230_2_R0_addr;
  wire  mem_230_2_R0_clk;
  wire [7:0] mem_230_2_R0_data;
  wire  mem_230_2_R0_en;
  wire [25:0] mem_230_2_W0_addr;
  wire  mem_230_2_W0_clk;
  wire [7:0] mem_230_2_W0_data;
  wire  mem_230_2_W0_en;
  wire  mem_230_2_W0_mask;
  wire [25:0] mem_230_3_R0_addr;
  wire  mem_230_3_R0_clk;
  wire [7:0] mem_230_3_R0_data;
  wire  mem_230_3_R0_en;
  wire [25:0] mem_230_3_W0_addr;
  wire  mem_230_3_W0_clk;
  wire [7:0] mem_230_3_W0_data;
  wire  mem_230_3_W0_en;
  wire  mem_230_3_W0_mask;
  wire [25:0] mem_230_4_R0_addr;
  wire  mem_230_4_R0_clk;
  wire [7:0] mem_230_4_R0_data;
  wire  mem_230_4_R0_en;
  wire [25:0] mem_230_4_W0_addr;
  wire  mem_230_4_W0_clk;
  wire [7:0] mem_230_4_W0_data;
  wire  mem_230_4_W0_en;
  wire  mem_230_4_W0_mask;
  wire [25:0] mem_230_5_R0_addr;
  wire  mem_230_5_R0_clk;
  wire [7:0] mem_230_5_R0_data;
  wire  mem_230_5_R0_en;
  wire [25:0] mem_230_5_W0_addr;
  wire  mem_230_5_W0_clk;
  wire [7:0] mem_230_5_W0_data;
  wire  mem_230_5_W0_en;
  wire  mem_230_5_W0_mask;
  wire [25:0] mem_230_6_R0_addr;
  wire  mem_230_6_R0_clk;
  wire [7:0] mem_230_6_R0_data;
  wire  mem_230_6_R0_en;
  wire [25:0] mem_230_6_W0_addr;
  wire  mem_230_6_W0_clk;
  wire [7:0] mem_230_6_W0_data;
  wire  mem_230_6_W0_en;
  wire  mem_230_6_W0_mask;
  wire [25:0] mem_230_7_R0_addr;
  wire  mem_230_7_R0_clk;
  wire [7:0] mem_230_7_R0_data;
  wire  mem_230_7_R0_en;
  wire [25:0] mem_230_7_W0_addr;
  wire  mem_230_7_W0_clk;
  wire [7:0] mem_230_7_W0_data;
  wire  mem_230_7_W0_en;
  wire  mem_230_7_W0_mask;
  wire [25:0] mem_231_0_R0_addr;
  wire  mem_231_0_R0_clk;
  wire [7:0] mem_231_0_R0_data;
  wire  mem_231_0_R0_en;
  wire [25:0] mem_231_0_W0_addr;
  wire  mem_231_0_W0_clk;
  wire [7:0] mem_231_0_W0_data;
  wire  mem_231_0_W0_en;
  wire  mem_231_0_W0_mask;
  wire [25:0] mem_231_1_R0_addr;
  wire  mem_231_1_R0_clk;
  wire [7:0] mem_231_1_R0_data;
  wire  mem_231_1_R0_en;
  wire [25:0] mem_231_1_W0_addr;
  wire  mem_231_1_W0_clk;
  wire [7:0] mem_231_1_W0_data;
  wire  mem_231_1_W0_en;
  wire  mem_231_1_W0_mask;
  wire [25:0] mem_231_2_R0_addr;
  wire  mem_231_2_R0_clk;
  wire [7:0] mem_231_2_R0_data;
  wire  mem_231_2_R0_en;
  wire [25:0] mem_231_2_W0_addr;
  wire  mem_231_2_W0_clk;
  wire [7:0] mem_231_2_W0_data;
  wire  mem_231_2_W0_en;
  wire  mem_231_2_W0_mask;
  wire [25:0] mem_231_3_R0_addr;
  wire  mem_231_3_R0_clk;
  wire [7:0] mem_231_3_R0_data;
  wire  mem_231_3_R0_en;
  wire [25:0] mem_231_3_W0_addr;
  wire  mem_231_3_W0_clk;
  wire [7:0] mem_231_3_W0_data;
  wire  mem_231_3_W0_en;
  wire  mem_231_3_W0_mask;
  wire [25:0] mem_231_4_R0_addr;
  wire  mem_231_4_R0_clk;
  wire [7:0] mem_231_4_R0_data;
  wire  mem_231_4_R0_en;
  wire [25:0] mem_231_4_W0_addr;
  wire  mem_231_4_W0_clk;
  wire [7:0] mem_231_4_W0_data;
  wire  mem_231_4_W0_en;
  wire  mem_231_4_W0_mask;
  wire [25:0] mem_231_5_R0_addr;
  wire  mem_231_5_R0_clk;
  wire [7:0] mem_231_5_R0_data;
  wire  mem_231_5_R0_en;
  wire [25:0] mem_231_5_W0_addr;
  wire  mem_231_5_W0_clk;
  wire [7:0] mem_231_5_W0_data;
  wire  mem_231_5_W0_en;
  wire  mem_231_5_W0_mask;
  wire [25:0] mem_231_6_R0_addr;
  wire  mem_231_6_R0_clk;
  wire [7:0] mem_231_6_R0_data;
  wire  mem_231_6_R0_en;
  wire [25:0] mem_231_6_W0_addr;
  wire  mem_231_6_W0_clk;
  wire [7:0] mem_231_6_W0_data;
  wire  mem_231_6_W0_en;
  wire  mem_231_6_W0_mask;
  wire [25:0] mem_231_7_R0_addr;
  wire  mem_231_7_R0_clk;
  wire [7:0] mem_231_7_R0_data;
  wire  mem_231_7_R0_en;
  wire [25:0] mem_231_7_W0_addr;
  wire  mem_231_7_W0_clk;
  wire [7:0] mem_231_7_W0_data;
  wire  mem_231_7_W0_en;
  wire  mem_231_7_W0_mask;
  wire [25:0] mem_232_0_R0_addr;
  wire  mem_232_0_R0_clk;
  wire [7:0] mem_232_0_R0_data;
  wire  mem_232_0_R0_en;
  wire [25:0] mem_232_0_W0_addr;
  wire  mem_232_0_W0_clk;
  wire [7:0] mem_232_0_W0_data;
  wire  mem_232_0_W0_en;
  wire  mem_232_0_W0_mask;
  wire [25:0] mem_232_1_R0_addr;
  wire  mem_232_1_R0_clk;
  wire [7:0] mem_232_1_R0_data;
  wire  mem_232_1_R0_en;
  wire [25:0] mem_232_1_W0_addr;
  wire  mem_232_1_W0_clk;
  wire [7:0] mem_232_1_W0_data;
  wire  mem_232_1_W0_en;
  wire  mem_232_1_W0_mask;
  wire [25:0] mem_232_2_R0_addr;
  wire  mem_232_2_R0_clk;
  wire [7:0] mem_232_2_R0_data;
  wire  mem_232_2_R0_en;
  wire [25:0] mem_232_2_W0_addr;
  wire  mem_232_2_W0_clk;
  wire [7:0] mem_232_2_W0_data;
  wire  mem_232_2_W0_en;
  wire  mem_232_2_W0_mask;
  wire [25:0] mem_232_3_R0_addr;
  wire  mem_232_3_R0_clk;
  wire [7:0] mem_232_3_R0_data;
  wire  mem_232_3_R0_en;
  wire [25:0] mem_232_3_W0_addr;
  wire  mem_232_3_W0_clk;
  wire [7:0] mem_232_3_W0_data;
  wire  mem_232_3_W0_en;
  wire  mem_232_3_W0_mask;
  wire [25:0] mem_232_4_R0_addr;
  wire  mem_232_4_R0_clk;
  wire [7:0] mem_232_4_R0_data;
  wire  mem_232_4_R0_en;
  wire [25:0] mem_232_4_W0_addr;
  wire  mem_232_4_W0_clk;
  wire [7:0] mem_232_4_W0_data;
  wire  mem_232_4_W0_en;
  wire  mem_232_4_W0_mask;
  wire [25:0] mem_232_5_R0_addr;
  wire  mem_232_5_R0_clk;
  wire [7:0] mem_232_5_R0_data;
  wire  mem_232_5_R0_en;
  wire [25:0] mem_232_5_W0_addr;
  wire  mem_232_5_W0_clk;
  wire [7:0] mem_232_5_W0_data;
  wire  mem_232_5_W0_en;
  wire  mem_232_5_W0_mask;
  wire [25:0] mem_232_6_R0_addr;
  wire  mem_232_6_R0_clk;
  wire [7:0] mem_232_6_R0_data;
  wire  mem_232_6_R0_en;
  wire [25:0] mem_232_6_W0_addr;
  wire  mem_232_6_W0_clk;
  wire [7:0] mem_232_6_W0_data;
  wire  mem_232_6_W0_en;
  wire  mem_232_6_W0_mask;
  wire [25:0] mem_232_7_R0_addr;
  wire  mem_232_7_R0_clk;
  wire [7:0] mem_232_7_R0_data;
  wire  mem_232_7_R0_en;
  wire [25:0] mem_232_7_W0_addr;
  wire  mem_232_7_W0_clk;
  wire [7:0] mem_232_7_W0_data;
  wire  mem_232_7_W0_en;
  wire  mem_232_7_W0_mask;
  wire [25:0] mem_233_0_R0_addr;
  wire  mem_233_0_R0_clk;
  wire [7:0] mem_233_0_R0_data;
  wire  mem_233_0_R0_en;
  wire [25:0] mem_233_0_W0_addr;
  wire  mem_233_0_W0_clk;
  wire [7:0] mem_233_0_W0_data;
  wire  mem_233_0_W0_en;
  wire  mem_233_0_W0_mask;
  wire [25:0] mem_233_1_R0_addr;
  wire  mem_233_1_R0_clk;
  wire [7:0] mem_233_1_R0_data;
  wire  mem_233_1_R0_en;
  wire [25:0] mem_233_1_W0_addr;
  wire  mem_233_1_W0_clk;
  wire [7:0] mem_233_1_W0_data;
  wire  mem_233_1_W0_en;
  wire  mem_233_1_W0_mask;
  wire [25:0] mem_233_2_R0_addr;
  wire  mem_233_2_R0_clk;
  wire [7:0] mem_233_2_R0_data;
  wire  mem_233_2_R0_en;
  wire [25:0] mem_233_2_W0_addr;
  wire  mem_233_2_W0_clk;
  wire [7:0] mem_233_2_W0_data;
  wire  mem_233_2_W0_en;
  wire  mem_233_2_W0_mask;
  wire [25:0] mem_233_3_R0_addr;
  wire  mem_233_3_R0_clk;
  wire [7:0] mem_233_3_R0_data;
  wire  mem_233_3_R0_en;
  wire [25:0] mem_233_3_W0_addr;
  wire  mem_233_3_W0_clk;
  wire [7:0] mem_233_3_W0_data;
  wire  mem_233_3_W0_en;
  wire  mem_233_3_W0_mask;
  wire [25:0] mem_233_4_R0_addr;
  wire  mem_233_4_R0_clk;
  wire [7:0] mem_233_4_R0_data;
  wire  mem_233_4_R0_en;
  wire [25:0] mem_233_4_W0_addr;
  wire  mem_233_4_W0_clk;
  wire [7:0] mem_233_4_W0_data;
  wire  mem_233_4_W0_en;
  wire  mem_233_4_W0_mask;
  wire [25:0] mem_233_5_R0_addr;
  wire  mem_233_5_R0_clk;
  wire [7:0] mem_233_5_R0_data;
  wire  mem_233_5_R0_en;
  wire [25:0] mem_233_5_W0_addr;
  wire  mem_233_5_W0_clk;
  wire [7:0] mem_233_5_W0_data;
  wire  mem_233_5_W0_en;
  wire  mem_233_5_W0_mask;
  wire [25:0] mem_233_6_R0_addr;
  wire  mem_233_6_R0_clk;
  wire [7:0] mem_233_6_R0_data;
  wire  mem_233_6_R0_en;
  wire [25:0] mem_233_6_W0_addr;
  wire  mem_233_6_W0_clk;
  wire [7:0] mem_233_6_W0_data;
  wire  mem_233_6_W0_en;
  wire  mem_233_6_W0_mask;
  wire [25:0] mem_233_7_R0_addr;
  wire  mem_233_7_R0_clk;
  wire [7:0] mem_233_7_R0_data;
  wire  mem_233_7_R0_en;
  wire [25:0] mem_233_7_W0_addr;
  wire  mem_233_7_W0_clk;
  wire [7:0] mem_233_7_W0_data;
  wire  mem_233_7_W0_en;
  wire  mem_233_7_W0_mask;
  wire [25:0] mem_234_0_R0_addr;
  wire  mem_234_0_R0_clk;
  wire [7:0] mem_234_0_R0_data;
  wire  mem_234_0_R0_en;
  wire [25:0] mem_234_0_W0_addr;
  wire  mem_234_0_W0_clk;
  wire [7:0] mem_234_0_W0_data;
  wire  mem_234_0_W0_en;
  wire  mem_234_0_W0_mask;
  wire [25:0] mem_234_1_R0_addr;
  wire  mem_234_1_R0_clk;
  wire [7:0] mem_234_1_R0_data;
  wire  mem_234_1_R0_en;
  wire [25:0] mem_234_1_W0_addr;
  wire  mem_234_1_W0_clk;
  wire [7:0] mem_234_1_W0_data;
  wire  mem_234_1_W0_en;
  wire  mem_234_1_W0_mask;
  wire [25:0] mem_234_2_R0_addr;
  wire  mem_234_2_R0_clk;
  wire [7:0] mem_234_2_R0_data;
  wire  mem_234_2_R0_en;
  wire [25:0] mem_234_2_W0_addr;
  wire  mem_234_2_W0_clk;
  wire [7:0] mem_234_2_W0_data;
  wire  mem_234_2_W0_en;
  wire  mem_234_2_W0_mask;
  wire [25:0] mem_234_3_R0_addr;
  wire  mem_234_3_R0_clk;
  wire [7:0] mem_234_3_R0_data;
  wire  mem_234_3_R0_en;
  wire [25:0] mem_234_3_W0_addr;
  wire  mem_234_3_W0_clk;
  wire [7:0] mem_234_3_W0_data;
  wire  mem_234_3_W0_en;
  wire  mem_234_3_W0_mask;
  wire [25:0] mem_234_4_R0_addr;
  wire  mem_234_4_R0_clk;
  wire [7:0] mem_234_4_R0_data;
  wire  mem_234_4_R0_en;
  wire [25:0] mem_234_4_W0_addr;
  wire  mem_234_4_W0_clk;
  wire [7:0] mem_234_4_W0_data;
  wire  mem_234_4_W0_en;
  wire  mem_234_4_W0_mask;
  wire [25:0] mem_234_5_R0_addr;
  wire  mem_234_5_R0_clk;
  wire [7:0] mem_234_5_R0_data;
  wire  mem_234_5_R0_en;
  wire [25:0] mem_234_5_W0_addr;
  wire  mem_234_5_W0_clk;
  wire [7:0] mem_234_5_W0_data;
  wire  mem_234_5_W0_en;
  wire  mem_234_5_W0_mask;
  wire [25:0] mem_234_6_R0_addr;
  wire  mem_234_6_R0_clk;
  wire [7:0] mem_234_6_R0_data;
  wire  mem_234_6_R0_en;
  wire [25:0] mem_234_6_W0_addr;
  wire  mem_234_6_W0_clk;
  wire [7:0] mem_234_6_W0_data;
  wire  mem_234_6_W0_en;
  wire  mem_234_6_W0_mask;
  wire [25:0] mem_234_7_R0_addr;
  wire  mem_234_7_R0_clk;
  wire [7:0] mem_234_7_R0_data;
  wire  mem_234_7_R0_en;
  wire [25:0] mem_234_7_W0_addr;
  wire  mem_234_7_W0_clk;
  wire [7:0] mem_234_7_W0_data;
  wire  mem_234_7_W0_en;
  wire  mem_234_7_W0_mask;
  wire [25:0] mem_235_0_R0_addr;
  wire  mem_235_0_R0_clk;
  wire [7:0] mem_235_0_R0_data;
  wire  mem_235_0_R0_en;
  wire [25:0] mem_235_0_W0_addr;
  wire  mem_235_0_W0_clk;
  wire [7:0] mem_235_0_W0_data;
  wire  mem_235_0_W0_en;
  wire  mem_235_0_W0_mask;
  wire [25:0] mem_235_1_R0_addr;
  wire  mem_235_1_R0_clk;
  wire [7:0] mem_235_1_R0_data;
  wire  mem_235_1_R0_en;
  wire [25:0] mem_235_1_W0_addr;
  wire  mem_235_1_W0_clk;
  wire [7:0] mem_235_1_W0_data;
  wire  mem_235_1_W0_en;
  wire  mem_235_1_W0_mask;
  wire [25:0] mem_235_2_R0_addr;
  wire  mem_235_2_R0_clk;
  wire [7:0] mem_235_2_R0_data;
  wire  mem_235_2_R0_en;
  wire [25:0] mem_235_2_W0_addr;
  wire  mem_235_2_W0_clk;
  wire [7:0] mem_235_2_W0_data;
  wire  mem_235_2_W0_en;
  wire  mem_235_2_W0_mask;
  wire [25:0] mem_235_3_R0_addr;
  wire  mem_235_3_R0_clk;
  wire [7:0] mem_235_3_R0_data;
  wire  mem_235_3_R0_en;
  wire [25:0] mem_235_3_W0_addr;
  wire  mem_235_3_W0_clk;
  wire [7:0] mem_235_3_W0_data;
  wire  mem_235_3_W0_en;
  wire  mem_235_3_W0_mask;
  wire [25:0] mem_235_4_R0_addr;
  wire  mem_235_4_R0_clk;
  wire [7:0] mem_235_4_R0_data;
  wire  mem_235_4_R0_en;
  wire [25:0] mem_235_4_W0_addr;
  wire  mem_235_4_W0_clk;
  wire [7:0] mem_235_4_W0_data;
  wire  mem_235_4_W0_en;
  wire  mem_235_4_W0_mask;
  wire [25:0] mem_235_5_R0_addr;
  wire  mem_235_5_R0_clk;
  wire [7:0] mem_235_5_R0_data;
  wire  mem_235_5_R0_en;
  wire [25:0] mem_235_5_W0_addr;
  wire  mem_235_5_W0_clk;
  wire [7:0] mem_235_5_W0_data;
  wire  mem_235_5_W0_en;
  wire  mem_235_5_W0_mask;
  wire [25:0] mem_235_6_R0_addr;
  wire  mem_235_6_R0_clk;
  wire [7:0] mem_235_6_R0_data;
  wire  mem_235_6_R0_en;
  wire [25:0] mem_235_6_W0_addr;
  wire  mem_235_6_W0_clk;
  wire [7:0] mem_235_6_W0_data;
  wire  mem_235_6_W0_en;
  wire  mem_235_6_W0_mask;
  wire [25:0] mem_235_7_R0_addr;
  wire  mem_235_7_R0_clk;
  wire [7:0] mem_235_7_R0_data;
  wire  mem_235_7_R0_en;
  wire [25:0] mem_235_7_W0_addr;
  wire  mem_235_7_W0_clk;
  wire [7:0] mem_235_7_W0_data;
  wire  mem_235_7_W0_en;
  wire  mem_235_7_W0_mask;
  wire [25:0] mem_236_0_R0_addr;
  wire  mem_236_0_R0_clk;
  wire [7:0] mem_236_0_R0_data;
  wire  mem_236_0_R0_en;
  wire [25:0] mem_236_0_W0_addr;
  wire  mem_236_0_W0_clk;
  wire [7:0] mem_236_0_W0_data;
  wire  mem_236_0_W0_en;
  wire  mem_236_0_W0_mask;
  wire [25:0] mem_236_1_R0_addr;
  wire  mem_236_1_R0_clk;
  wire [7:0] mem_236_1_R0_data;
  wire  mem_236_1_R0_en;
  wire [25:0] mem_236_1_W0_addr;
  wire  mem_236_1_W0_clk;
  wire [7:0] mem_236_1_W0_data;
  wire  mem_236_1_W0_en;
  wire  mem_236_1_W0_mask;
  wire [25:0] mem_236_2_R0_addr;
  wire  mem_236_2_R0_clk;
  wire [7:0] mem_236_2_R0_data;
  wire  mem_236_2_R0_en;
  wire [25:0] mem_236_2_W0_addr;
  wire  mem_236_2_W0_clk;
  wire [7:0] mem_236_2_W0_data;
  wire  mem_236_2_W0_en;
  wire  mem_236_2_W0_mask;
  wire [25:0] mem_236_3_R0_addr;
  wire  mem_236_3_R0_clk;
  wire [7:0] mem_236_3_R0_data;
  wire  mem_236_3_R0_en;
  wire [25:0] mem_236_3_W0_addr;
  wire  mem_236_3_W0_clk;
  wire [7:0] mem_236_3_W0_data;
  wire  mem_236_3_W0_en;
  wire  mem_236_3_W0_mask;
  wire [25:0] mem_236_4_R0_addr;
  wire  mem_236_4_R0_clk;
  wire [7:0] mem_236_4_R0_data;
  wire  mem_236_4_R0_en;
  wire [25:0] mem_236_4_W0_addr;
  wire  mem_236_4_W0_clk;
  wire [7:0] mem_236_4_W0_data;
  wire  mem_236_4_W0_en;
  wire  mem_236_4_W0_mask;
  wire [25:0] mem_236_5_R0_addr;
  wire  mem_236_5_R0_clk;
  wire [7:0] mem_236_5_R0_data;
  wire  mem_236_5_R0_en;
  wire [25:0] mem_236_5_W0_addr;
  wire  mem_236_5_W0_clk;
  wire [7:0] mem_236_5_W0_data;
  wire  mem_236_5_W0_en;
  wire  mem_236_5_W0_mask;
  wire [25:0] mem_236_6_R0_addr;
  wire  mem_236_6_R0_clk;
  wire [7:0] mem_236_6_R0_data;
  wire  mem_236_6_R0_en;
  wire [25:0] mem_236_6_W0_addr;
  wire  mem_236_6_W0_clk;
  wire [7:0] mem_236_6_W0_data;
  wire  mem_236_6_W0_en;
  wire  mem_236_6_W0_mask;
  wire [25:0] mem_236_7_R0_addr;
  wire  mem_236_7_R0_clk;
  wire [7:0] mem_236_7_R0_data;
  wire  mem_236_7_R0_en;
  wire [25:0] mem_236_7_W0_addr;
  wire  mem_236_7_W0_clk;
  wire [7:0] mem_236_7_W0_data;
  wire  mem_236_7_W0_en;
  wire  mem_236_7_W0_mask;
  wire [25:0] mem_237_0_R0_addr;
  wire  mem_237_0_R0_clk;
  wire [7:0] mem_237_0_R0_data;
  wire  mem_237_0_R0_en;
  wire [25:0] mem_237_0_W0_addr;
  wire  mem_237_0_W0_clk;
  wire [7:0] mem_237_0_W0_data;
  wire  mem_237_0_W0_en;
  wire  mem_237_0_W0_mask;
  wire [25:0] mem_237_1_R0_addr;
  wire  mem_237_1_R0_clk;
  wire [7:0] mem_237_1_R0_data;
  wire  mem_237_1_R0_en;
  wire [25:0] mem_237_1_W0_addr;
  wire  mem_237_1_W0_clk;
  wire [7:0] mem_237_1_W0_data;
  wire  mem_237_1_W0_en;
  wire  mem_237_1_W0_mask;
  wire [25:0] mem_237_2_R0_addr;
  wire  mem_237_2_R0_clk;
  wire [7:0] mem_237_2_R0_data;
  wire  mem_237_2_R0_en;
  wire [25:0] mem_237_2_W0_addr;
  wire  mem_237_2_W0_clk;
  wire [7:0] mem_237_2_W0_data;
  wire  mem_237_2_W0_en;
  wire  mem_237_2_W0_mask;
  wire [25:0] mem_237_3_R0_addr;
  wire  mem_237_3_R0_clk;
  wire [7:0] mem_237_3_R0_data;
  wire  mem_237_3_R0_en;
  wire [25:0] mem_237_3_W0_addr;
  wire  mem_237_3_W0_clk;
  wire [7:0] mem_237_3_W0_data;
  wire  mem_237_3_W0_en;
  wire  mem_237_3_W0_mask;
  wire [25:0] mem_237_4_R0_addr;
  wire  mem_237_4_R0_clk;
  wire [7:0] mem_237_4_R0_data;
  wire  mem_237_4_R0_en;
  wire [25:0] mem_237_4_W0_addr;
  wire  mem_237_4_W0_clk;
  wire [7:0] mem_237_4_W0_data;
  wire  mem_237_4_W0_en;
  wire  mem_237_4_W0_mask;
  wire [25:0] mem_237_5_R0_addr;
  wire  mem_237_5_R0_clk;
  wire [7:0] mem_237_5_R0_data;
  wire  mem_237_5_R0_en;
  wire [25:0] mem_237_5_W0_addr;
  wire  mem_237_5_W0_clk;
  wire [7:0] mem_237_5_W0_data;
  wire  mem_237_5_W0_en;
  wire  mem_237_5_W0_mask;
  wire [25:0] mem_237_6_R0_addr;
  wire  mem_237_6_R0_clk;
  wire [7:0] mem_237_6_R0_data;
  wire  mem_237_6_R0_en;
  wire [25:0] mem_237_6_W0_addr;
  wire  mem_237_6_W0_clk;
  wire [7:0] mem_237_6_W0_data;
  wire  mem_237_6_W0_en;
  wire  mem_237_6_W0_mask;
  wire [25:0] mem_237_7_R0_addr;
  wire  mem_237_7_R0_clk;
  wire [7:0] mem_237_7_R0_data;
  wire  mem_237_7_R0_en;
  wire [25:0] mem_237_7_W0_addr;
  wire  mem_237_7_W0_clk;
  wire [7:0] mem_237_7_W0_data;
  wire  mem_237_7_W0_en;
  wire  mem_237_7_W0_mask;
  wire [25:0] mem_238_0_R0_addr;
  wire  mem_238_0_R0_clk;
  wire [7:0] mem_238_0_R0_data;
  wire  mem_238_0_R0_en;
  wire [25:0] mem_238_0_W0_addr;
  wire  mem_238_0_W0_clk;
  wire [7:0] mem_238_0_W0_data;
  wire  mem_238_0_W0_en;
  wire  mem_238_0_W0_mask;
  wire [25:0] mem_238_1_R0_addr;
  wire  mem_238_1_R0_clk;
  wire [7:0] mem_238_1_R0_data;
  wire  mem_238_1_R0_en;
  wire [25:0] mem_238_1_W0_addr;
  wire  mem_238_1_W0_clk;
  wire [7:0] mem_238_1_W0_data;
  wire  mem_238_1_W0_en;
  wire  mem_238_1_W0_mask;
  wire [25:0] mem_238_2_R0_addr;
  wire  mem_238_2_R0_clk;
  wire [7:0] mem_238_2_R0_data;
  wire  mem_238_2_R0_en;
  wire [25:0] mem_238_2_W0_addr;
  wire  mem_238_2_W0_clk;
  wire [7:0] mem_238_2_W0_data;
  wire  mem_238_2_W0_en;
  wire  mem_238_2_W0_mask;
  wire [25:0] mem_238_3_R0_addr;
  wire  mem_238_3_R0_clk;
  wire [7:0] mem_238_3_R0_data;
  wire  mem_238_3_R0_en;
  wire [25:0] mem_238_3_W0_addr;
  wire  mem_238_3_W0_clk;
  wire [7:0] mem_238_3_W0_data;
  wire  mem_238_3_W0_en;
  wire  mem_238_3_W0_mask;
  wire [25:0] mem_238_4_R0_addr;
  wire  mem_238_4_R0_clk;
  wire [7:0] mem_238_4_R0_data;
  wire  mem_238_4_R0_en;
  wire [25:0] mem_238_4_W0_addr;
  wire  mem_238_4_W0_clk;
  wire [7:0] mem_238_4_W0_data;
  wire  mem_238_4_W0_en;
  wire  mem_238_4_W0_mask;
  wire [25:0] mem_238_5_R0_addr;
  wire  mem_238_5_R0_clk;
  wire [7:0] mem_238_5_R0_data;
  wire  mem_238_5_R0_en;
  wire [25:0] mem_238_5_W0_addr;
  wire  mem_238_5_W0_clk;
  wire [7:0] mem_238_5_W0_data;
  wire  mem_238_5_W0_en;
  wire  mem_238_5_W0_mask;
  wire [25:0] mem_238_6_R0_addr;
  wire  mem_238_6_R0_clk;
  wire [7:0] mem_238_6_R0_data;
  wire  mem_238_6_R0_en;
  wire [25:0] mem_238_6_W0_addr;
  wire  mem_238_6_W0_clk;
  wire [7:0] mem_238_6_W0_data;
  wire  mem_238_6_W0_en;
  wire  mem_238_6_W0_mask;
  wire [25:0] mem_238_7_R0_addr;
  wire  mem_238_7_R0_clk;
  wire [7:0] mem_238_7_R0_data;
  wire  mem_238_7_R0_en;
  wire [25:0] mem_238_7_W0_addr;
  wire  mem_238_7_W0_clk;
  wire [7:0] mem_238_7_W0_data;
  wire  mem_238_7_W0_en;
  wire  mem_238_7_W0_mask;
  wire [25:0] mem_239_0_R0_addr;
  wire  mem_239_0_R0_clk;
  wire [7:0] mem_239_0_R0_data;
  wire  mem_239_0_R0_en;
  wire [25:0] mem_239_0_W0_addr;
  wire  mem_239_0_W0_clk;
  wire [7:0] mem_239_0_W0_data;
  wire  mem_239_0_W0_en;
  wire  mem_239_0_W0_mask;
  wire [25:0] mem_239_1_R0_addr;
  wire  mem_239_1_R0_clk;
  wire [7:0] mem_239_1_R0_data;
  wire  mem_239_1_R0_en;
  wire [25:0] mem_239_1_W0_addr;
  wire  mem_239_1_W0_clk;
  wire [7:0] mem_239_1_W0_data;
  wire  mem_239_1_W0_en;
  wire  mem_239_1_W0_mask;
  wire [25:0] mem_239_2_R0_addr;
  wire  mem_239_2_R0_clk;
  wire [7:0] mem_239_2_R0_data;
  wire  mem_239_2_R0_en;
  wire [25:0] mem_239_2_W0_addr;
  wire  mem_239_2_W0_clk;
  wire [7:0] mem_239_2_W0_data;
  wire  mem_239_2_W0_en;
  wire  mem_239_2_W0_mask;
  wire [25:0] mem_239_3_R0_addr;
  wire  mem_239_3_R0_clk;
  wire [7:0] mem_239_3_R0_data;
  wire  mem_239_3_R0_en;
  wire [25:0] mem_239_3_W0_addr;
  wire  mem_239_3_W0_clk;
  wire [7:0] mem_239_3_W0_data;
  wire  mem_239_3_W0_en;
  wire  mem_239_3_W0_mask;
  wire [25:0] mem_239_4_R0_addr;
  wire  mem_239_4_R0_clk;
  wire [7:0] mem_239_4_R0_data;
  wire  mem_239_4_R0_en;
  wire [25:0] mem_239_4_W0_addr;
  wire  mem_239_4_W0_clk;
  wire [7:0] mem_239_4_W0_data;
  wire  mem_239_4_W0_en;
  wire  mem_239_4_W0_mask;
  wire [25:0] mem_239_5_R0_addr;
  wire  mem_239_5_R0_clk;
  wire [7:0] mem_239_5_R0_data;
  wire  mem_239_5_R0_en;
  wire [25:0] mem_239_5_W0_addr;
  wire  mem_239_5_W0_clk;
  wire [7:0] mem_239_5_W0_data;
  wire  mem_239_5_W0_en;
  wire  mem_239_5_W0_mask;
  wire [25:0] mem_239_6_R0_addr;
  wire  mem_239_6_R0_clk;
  wire [7:0] mem_239_6_R0_data;
  wire  mem_239_6_R0_en;
  wire [25:0] mem_239_6_W0_addr;
  wire  mem_239_6_W0_clk;
  wire [7:0] mem_239_6_W0_data;
  wire  mem_239_6_W0_en;
  wire  mem_239_6_W0_mask;
  wire [25:0] mem_239_7_R0_addr;
  wire  mem_239_7_R0_clk;
  wire [7:0] mem_239_7_R0_data;
  wire  mem_239_7_R0_en;
  wire [25:0] mem_239_7_W0_addr;
  wire  mem_239_7_W0_clk;
  wire [7:0] mem_239_7_W0_data;
  wire  mem_239_7_W0_en;
  wire  mem_239_7_W0_mask;
  wire [25:0] mem_240_0_R0_addr;
  wire  mem_240_0_R0_clk;
  wire [7:0] mem_240_0_R0_data;
  wire  mem_240_0_R0_en;
  wire [25:0] mem_240_0_W0_addr;
  wire  mem_240_0_W0_clk;
  wire [7:0] mem_240_0_W0_data;
  wire  mem_240_0_W0_en;
  wire  mem_240_0_W0_mask;
  wire [25:0] mem_240_1_R0_addr;
  wire  mem_240_1_R0_clk;
  wire [7:0] mem_240_1_R0_data;
  wire  mem_240_1_R0_en;
  wire [25:0] mem_240_1_W0_addr;
  wire  mem_240_1_W0_clk;
  wire [7:0] mem_240_1_W0_data;
  wire  mem_240_1_W0_en;
  wire  mem_240_1_W0_mask;
  wire [25:0] mem_240_2_R0_addr;
  wire  mem_240_2_R0_clk;
  wire [7:0] mem_240_2_R0_data;
  wire  mem_240_2_R0_en;
  wire [25:0] mem_240_2_W0_addr;
  wire  mem_240_2_W0_clk;
  wire [7:0] mem_240_2_W0_data;
  wire  mem_240_2_W0_en;
  wire  mem_240_2_W0_mask;
  wire [25:0] mem_240_3_R0_addr;
  wire  mem_240_3_R0_clk;
  wire [7:0] mem_240_3_R0_data;
  wire  mem_240_3_R0_en;
  wire [25:0] mem_240_3_W0_addr;
  wire  mem_240_3_W0_clk;
  wire [7:0] mem_240_3_W0_data;
  wire  mem_240_3_W0_en;
  wire  mem_240_3_W0_mask;
  wire [25:0] mem_240_4_R0_addr;
  wire  mem_240_4_R0_clk;
  wire [7:0] mem_240_4_R0_data;
  wire  mem_240_4_R0_en;
  wire [25:0] mem_240_4_W0_addr;
  wire  mem_240_4_W0_clk;
  wire [7:0] mem_240_4_W0_data;
  wire  mem_240_4_W0_en;
  wire  mem_240_4_W0_mask;
  wire [25:0] mem_240_5_R0_addr;
  wire  mem_240_5_R0_clk;
  wire [7:0] mem_240_5_R0_data;
  wire  mem_240_5_R0_en;
  wire [25:0] mem_240_5_W0_addr;
  wire  mem_240_5_W0_clk;
  wire [7:0] mem_240_5_W0_data;
  wire  mem_240_5_W0_en;
  wire  mem_240_5_W0_mask;
  wire [25:0] mem_240_6_R0_addr;
  wire  mem_240_6_R0_clk;
  wire [7:0] mem_240_6_R0_data;
  wire  mem_240_6_R0_en;
  wire [25:0] mem_240_6_W0_addr;
  wire  mem_240_6_W0_clk;
  wire [7:0] mem_240_6_W0_data;
  wire  mem_240_6_W0_en;
  wire  mem_240_6_W0_mask;
  wire [25:0] mem_240_7_R0_addr;
  wire  mem_240_7_R0_clk;
  wire [7:0] mem_240_7_R0_data;
  wire  mem_240_7_R0_en;
  wire [25:0] mem_240_7_W0_addr;
  wire  mem_240_7_W0_clk;
  wire [7:0] mem_240_7_W0_data;
  wire  mem_240_7_W0_en;
  wire  mem_240_7_W0_mask;
  wire [25:0] mem_241_0_R0_addr;
  wire  mem_241_0_R0_clk;
  wire [7:0] mem_241_0_R0_data;
  wire  mem_241_0_R0_en;
  wire [25:0] mem_241_0_W0_addr;
  wire  mem_241_0_W0_clk;
  wire [7:0] mem_241_0_W0_data;
  wire  mem_241_0_W0_en;
  wire  mem_241_0_W0_mask;
  wire [25:0] mem_241_1_R0_addr;
  wire  mem_241_1_R0_clk;
  wire [7:0] mem_241_1_R0_data;
  wire  mem_241_1_R0_en;
  wire [25:0] mem_241_1_W0_addr;
  wire  mem_241_1_W0_clk;
  wire [7:0] mem_241_1_W0_data;
  wire  mem_241_1_W0_en;
  wire  mem_241_1_W0_mask;
  wire [25:0] mem_241_2_R0_addr;
  wire  mem_241_2_R0_clk;
  wire [7:0] mem_241_2_R0_data;
  wire  mem_241_2_R0_en;
  wire [25:0] mem_241_2_W0_addr;
  wire  mem_241_2_W0_clk;
  wire [7:0] mem_241_2_W0_data;
  wire  mem_241_2_W0_en;
  wire  mem_241_2_W0_mask;
  wire [25:0] mem_241_3_R0_addr;
  wire  mem_241_3_R0_clk;
  wire [7:0] mem_241_3_R0_data;
  wire  mem_241_3_R0_en;
  wire [25:0] mem_241_3_W0_addr;
  wire  mem_241_3_W0_clk;
  wire [7:0] mem_241_3_W0_data;
  wire  mem_241_3_W0_en;
  wire  mem_241_3_W0_mask;
  wire [25:0] mem_241_4_R0_addr;
  wire  mem_241_4_R0_clk;
  wire [7:0] mem_241_4_R0_data;
  wire  mem_241_4_R0_en;
  wire [25:0] mem_241_4_W0_addr;
  wire  mem_241_4_W0_clk;
  wire [7:0] mem_241_4_W0_data;
  wire  mem_241_4_W0_en;
  wire  mem_241_4_W0_mask;
  wire [25:0] mem_241_5_R0_addr;
  wire  mem_241_5_R0_clk;
  wire [7:0] mem_241_5_R0_data;
  wire  mem_241_5_R0_en;
  wire [25:0] mem_241_5_W0_addr;
  wire  mem_241_5_W0_clk;
  wire [7:0] mem_241_5_W0_data;
  wire  mem_241_5_W0_en;
  wire  mem_241_5_W0_mask;
  wire [25:0] mem_241_6_R0_addr;
  wire  mem_241_6_R0_clk;
  wire [7:0] mem_241_6_R0_data;
  wire  mem_241_6_R0_en;
  wire [25:0] mem_241_6_W0_addr;
  wire  mem_241_6_W0_clk;
  wire [7:0] mem_241_6_W0_data;
  wire  mem_241_6_W0_en;
  wire  mem_241_6_W0_mask;
  wire [25:0] mem_241_7_R0_addr;
  wire  mem_241_7_R0_clk;
  wire [7:0] mem_241_7_R0_data;
  wire  mem_241_7_R0_en;
  wire [25:0] mem_241_7_W0_addr;
  wire  mem_241_7_W0_clk;
  wire [7:0] mem_241_7_W0_data;
  wire  mem_241_7_W0_en;
  wire  mem_241_7_W0_mask;
  wire [25:0] mem_242_0_R0_addr;
  wire  mem_242_0_R0_clk;
  wire [7:0] mem_242_0_R0_data;
  wire  mem_242_0_R0_en;
  wire [25:0] mem_242_0_W0_addr;
  wire  mem_242_0_W0_clk;
  wire [7:0] mem_242_0_W0_data;
  wire  mem_242_0_W0_en;
  wire  mem_242_0_W0_mask;
  wire [25:0] mem_242_1_R0_addr;
  wire  mem_242_1_R0_clk;
  wire [7:0] mem_242_1_R0_data;
  wire  mem_242_1_R0_en;
  wire [25:0] mem_242_1_W0_addr;
  wire  mem_242_1_W0_clk;
  wire [7:0] mem_242_1_W0_data;
  wire  mem_242_1_W0_en;
  wire  mem_242_1_W0_mask;
  wire [25:0] mem_242_2_R0_addr;
  wire  mem_242_2_R0_clk;
  wire [7:0] mem_242_2_R0_data;
  wire  mem_242_2_R0_en;
  wire [25:0] mem_242_2_W0_addr;
  wire  mem_242_2_W0_clk;
  wire [7:0] mem_242_2_W0_data;
  wire  mem_242_2_W0_en;
  wire  mem_242_2_W0_mask;
  wire [25:0] mem_242_3_R0_addr;
  wire  mem_242_3_R0_clk;
  wire [7:0] mem_242_3_R0_data;
  wire  mem_242_3_R0_en;
  wire [25:0] mem_242_3_W0_addr;
  wire  mem_242_3_W0_clk;
  wire [7:0] mem_242_3_W0_data;
  wire  mem_242_3_W0_en;
  wire  mem_242_3_W0_mask;
  wire [25:0] mem_242_4_R0_addr;
  wire  mem_242_4_R0_clk;
  wire [7:0] mem_242_4_R0_data;
  wire  mem_242_4_R0_en;
  wire [25:0] mem_242_4_W0_addr;
  wire  mem_242_4_W0_clk;
  wire [7:0] mem_242_4_W0_data;
  wire  mem_242_4_W0_en;
  wire  mem_242_4_W0_mask;
  wire [25:0] mem_242_5_R0_addr;
  wire  mem_242_5_R0_clk;
  wire [7:0] mem_242_5_R0_data;
  wire  mem_242_5_R0_en;
  wire [25:0] mem_242_5_W0_addr;
  wire  mem_242_5_W0_clk;
  wire [7:0] mem_242_5_W0_data;
  wire  mem_242_5_W0_en;
  wire  mem_242_5_W0_mask;
  wire [25:0] mem_242_6_R0_addr;
  wire  mem_242_6_R0_clk;
  wire [7:0] mem_242_6_R0_data;
  wire  mem_242_6_R0_en;
  wire [25:0] mem_242_6_W0_addr;
  wire  mem_242_6_W0_clk;
  wire [7:0] mem_242_6_W0_data;
  wire  mem_242_6_W0_en;
  wire  mem_242_6_W0_mask;
  wire [25:0] mem_242_7_R0_addr;
  wire  mem_242_7_R0_clk;
  wire [7:0] mem_242_7_R0_data;
  wire  mem_242_7_R0_en;
  wire [25:0] mem_242_7_W0_addr;
  wire  mem_242_7_W0_clk;
  wire [7:0] mem_242_7_W0_data;
  wire  mem_242_7_W0_en;
  wire  mem_242_7_W0_mask;
  wire [25:0] mem_243_0_R0_addr;
  wire  mem_243_0_R0_clk;
  wire [7:0] mem_243_0_R0_data;
  wire  mem_243_0_R0_en;
  wire [25:0] mem_243_0_W0_addr;
  wire  mem_243_0_W0_clk;
  wire [7:0] mem_243_0_W0_data;
  wire  mem_243_0_W0_en;
  wire  mem_243_0_W0_mask;
  wire [25:0] mem_243_1_R0_addr;
  wire  mem_243_1_R0_clk;
  wire [7:0] mem_243_1_R0_data;
  wire  mem_243_1_R0_en;
  wire [25:0] mem_243_1_W0_addr;
  wire  mem_243_1_W0_clk;
  wire [7:0] mem_243_1_W0_data;
  wire  mem_243_1_W0_en;
  wire  mem_243_1_W0_mask;
  wire [25:0] mem_243_2_R0_addr;
  wire  mem_243_2_R0_clk;
  wire [7:0] mem_243_2_R0_data;
  wire  mem_243_2_R0_en;
  wire [25:0] mem_243_2_W0_addr;
  wire  mem_243_2_W0_clk;
  wire [7:0] mem_243_2_W0_data;
  wire  mem_243_2_W0_en;
  wire  mem_243_2_W0_mask;
  wire [25:0] mem_243_3_R0_addr;
  wire  mem_243_3_R0_clk;
  wire [7:0] mem_243_3_R0_data;
  wire  mem_243_3_R0_en;
  wire [25:0] mem_243_3_W0_addr;
  wire  mem_243_3_W0_clk;
  wire [7:0] mem_243_3_W0_data;
  wire  mem_243_3_W0_en;
  wire  mem_243_3_W0_mask;
  wire [25:0] mem_243_4_R0_addr;
  wire  mem_243_4_R0_clk;
  wire [7:0] mem_243_4_R0_data;
  wire  mem_243_4_R0_en;
  wire [25:0] mem_243_4_W0_addr;
  wire  mem_243_4_W0_clk;
  wire [7:0] mem_243_4_W0_data;
  wire  mem_243_4_W0_en;
  wire  mem_243_4_W0_mask;
  wire [25:0] mem_243_5_R0_addr;
  wire  mem_243_5_R0_clk;
  wire [7:0] mem_243_5_R0_data;
  wire  mem_243_5_R0_en;
  wire [25:0] mem_243_5_W0_addr;
  wire  mem_243_5_W0_clk;
  wire [7:0] mem_243_5_W0_data;
  wire  mem_243_5_W0_en;
  wire  mem_243_5_W0_mask;
  wire [25:0] mem_243_6_R0_addr;
  wire  mem_243_6_R0_clk;
  wire [7:0] mem_243_6_R0_data;
  wire  mem_243_6_R0_en;
  wire [25:0] mem_243_6_W0_addr;
  wire  mem_243_6_W0_clk;
  wire [7:0] mem_243_6_W0_data;
  wire  mem_243_6_W0_en;
  wire  mem_243_6_W0_mask;
  wire [25:0] mem_243_7_R0_addr;
  wire  mem_243_7_R0_clk;
  wire [7:0] mem_243_7_R0_data;
  wire  mem_243_7_R0_en;
  wire [25:0] mem_243_7_W0_addr;
  wire  mem_243_7_W0_clk;
  wire [7:0] mem_243_7_W0_data;
  wire  mem_243_7_W0_en;
  wire  mem_243_7_W0_mask;
  wire [25:0] mem_244_0_R0_addr;
  wire  mem_244_0_R0_clk;
  wire [7:0] mem_244_0_R0_data;
  wire  mem_244_0_R0_en;
  wire [25:0] mem_244_0_W0_addr;
  wire  mem_244_0_W0_clk;
  wire [7:0] mem_244_0_W0_data;
  wire  mem_244_0_W0_en;
  wire  mem_244_0_W0_mask;
  wire [25:0] mem_244_1_R0_addr;
  wire  mem_244_1_R0_clk;
  wire [7:0] mem_244_1_R0_data;
  wire  mem_244_1_R0_en;
  wire [25:0] mem_244_1_W0_addr;
  wire  mem_244_1_W0_clk;
  wire [7:0] mem_244_1_W0_data;
  wire  mem_244_1_W0_en;
  wire  mem_244_1_W0_mask;
  wire [25:0] mem_244_2_R0_addr;
  wire  mem_244_2_R0_clk;
  wire [7:0] mem_244_2_R0_data;
  wire  mem_244_2_R0_en;
  wire [25:0] mem_244_2_W0_addr;
  wire  mem_244_2_W0_clk;
  wire [7:0] mem_244_2_W0_data;
  wire  mem_244_2_W0_en;
  wire  mem_244_2_W0_mask;
  wire [25:0] mem_244_3_R0_addr;
  wire  mem_244_3_R0_clk;
  wire [7:0] mem_244_3_R0_data;
  wire  mem_244_3_R0_en;
  wire [25:0] mem_244_3_W0_addr;
  wire  mem_244_3_W0_clk;
  wire [7:0] mem_244_3_W0_data;
  wire  mem_244_3_W0_en;
  wire  mem_244_3_W0_mask;
  wire [25:0] mem_244_4_R0_addr;
  wire  mem_244_4_R0_clk;
  wire [7:0] mem_244_4_R0_data;
  wire  mem_244_4_R0_en;
  wire [25:0] mem_244_4_W0_addr;
  wire  mem_244_4_W0_clk;
  wire [7:0] mem_244_4_W0_data;
  wire  mem_244_4_W0_en;
  wire  mem_244_4_W0_mask;
  wire [25:0] mem_244_5_R0_addr;
  wire  mem_244_5_R0_clk;
  wire [7:0] mem_244_5_R0_data;
  wire  mem_244_5_R0_en;
  wire [25:0] mem_244_5_W0_addr;
  wire  mem_244_5_W0_clk;
  wire [7:0] mem_244_5_W0_data;
  wire  mem_244_5_W0_en;
  wire  mem_244_5_W0_mask;
  wire [25:0] mem_244_6_R0_addr;
  wire  mem_244_6_R0_clk;
  wire [7:0] mem_244_6_R0_data;
  wire  mem_244_6_R0_en;
  wire [25:0] mem_244_6_W0_addr;
  wire  mem_244_6_W0_clk;
  wire [7:0] mem_244_6_W0_data;
  wire  mem_244_6_W0_en;
  wire  mem_244_6_W0_mask;
  wire [25:0] mem_244_7_R0_addr;
  wire  mem_244_7_R0_clk;
  wire [7:0] mem_244_7_R0_data;
  wire  mem_244_7_R0_en;
  wire [25:0] mem_244_7_W0_addr;
  wire  mem_244_7_W0_clk;
  wire [7:0] mem_244_7_W0_data;
  wire  mem_244_7_W0_en;
  wire  mem_244_7_W0_mask;
  wire [25:0] mem_245_0_R0_addr;
  wire  mem_245_0_R0_clk;
  wire [7:0] mem_245_0_R0_data;
  wire  mem_245_0_R0_en;
  wire [25:0] mem_245_0_W0_addr;
  wire  mem_245_0_W0_clk;
  wire [7:0] mem_245_0_W0_data;
  wire  mem_245_0_W0_en;
  wire  mem_245_0_W0_mask;
  wire [25:0] mem_245_1_R0_addr;
  wire  mem_245_1_R0_clk;
  wire [7:0] mem_245_1_R0_data;
  wire  mem_245_1_R0_en;
  wire [25:0] mem_245_1_W0_addr;
  wire  mem_245_1_W0_clk;
  wire [7:0] mem_245_1_W0_data;
  wire  mem_245_1_W0_en;
  wire  mem_245_1_W0_mask;
  wire [25:0] mem_245_2_R0_addr;
  wire  mem_245_2_R0_clk;
  wire [7:0] mem_245_2_R0_data;
  wire  mem_245_2_R0_en;
  wire [25:0] mem_245_2_W0_addr;
  wire  mem_245_2_W0_clk;
  wire [7:0] mem_245_2_W0_data;
  wire  mem_245_2_W0_en;
  wire  mem_245_2_W0_mask;
  wire [25:0] mem_245_3_R0_addr;
  wire  mem_245_3_R0_clk;
  wire [7:0] mem_245_3_R0_data;
  wire  mem_245_3_R0_en;
  wire [25:0] mem_245_3_W0_addr;
  wire  mem_245_3_W0_clk;
  wire [7:0] mem_245_3_W0_data;
  wire  mem_245_3_W0_en;
  wire  mem_245_3_W0_mask;
  wire [25:0] mem_245_4_R0_addr;
  wire  mem_245_4_R0_clk;
  wire [7:0] mem_245_4_R0_data;
  wire  mem_245_4_R0_en;
  wire [25:0] mem_245_4_W0_addr;
  wire  mem_245_4_W0_clk;
  wire [7:0] mem_245_4_W0_data;
  wire  mem_245_4_W0_en;
  wire  mem_245_4_W0_mask;
  wire [25:0] mem_245_5_R0_addr;
  wire  mem_245_5_R0_clk;
  wire [7:0] mem_245_5_R0_data;
  wire  mem_245_5_R0_en;
  wire [25:0] mem_245_5_W0_addr;
  wire  mem_245_5_W0_clk;
  wire [7:0] mem_245_5_W0_data;
  wire  mem_245_5_W0_en;
  wire  mem_245_5_W0_mask;
  wire [25:0] mem_245_6_R0_addr;
  wire  mem_245_6_R0_clk;
  wire [7:0] mem_245_6_R0_data;
  wire  mem_245_6_R0_en;
  wire [25:0] mem_245_6_W0_addr;
  wire  mem_245_6_W0_clk;
  wire [7:0] mem_245_6_W0_data;
  wire  mem_245_6_W0_en;
  wire  mem_245_6_W0_mask;
  wire [25:0] mem_245_7_R0_addr;
  wire  mem_245_7_R0_clk;
  wire [7:0] mem_245_7_R0_data;
  wire  mem_245_7_R0_en;
  wire [25:0] mem_245_7_W0_addr;
  wire  mem_245_7_W0_clk;
  wire [7:0] mem_245_7_W0_data;
  wire  mem_245_7_W0_en;
  wire  mem_245_7_W0_mask;
  wire [25:0] mem_246_0_R0_addr;
  wire  mem_246_0_R0_clk;
  wire [7:0] mem_246_0_R0_data;
  wire  mem_246_0_R0_en;
  wire [25:0] mem_246_0_W0_addr;
  wire  mem_246_0_W0_clk;
  wire [7:0] mem_246_0_W0_data;
  wire  mem_246_0_W0_en;
  wire  mem_246_0_W0_mask;
  wire [25:0] mem_246_1_R0_addr;
  wire  mem_246_1_R0_clk;
  wire [7:0] mem_246_1_R0_data;
  wire  mem_246_1_R0_en;
  wire [25:0] mem_246_1_W0_addr;
  wire  mem_246_1_W0_clk;
  wire [7:0] mem_246_1_W0_data;
  wire  mem_246_1_W0_en;
  wire  mem_246_1_W0_mask;
  wire [25:0] mem_246_2_R0_addr;
  wire  mem_246_2_R0_clk;
  wire [7:0] mem_246_2_R0_data;
  wire  mem_246_2_R0_en;
  wire [25:0] mem_246_2_W0_addr;
  wire  mem_246_2_W0_clk;
  wire [7:0] mem_246_2_W0_data;
  wire  mem_246_2_W0_en;
  wire  mem_246_2_W0_mask;
  wire [25:0] mem_246_3_R0_addr;
  wire  mem_246_3_R0_clk;
  wire [7:0] mem_246_3_R0_data;
  wire  mem_246_3_R0_en;
  wire [25:0] mem_246_3_W0_addr;
  wire  mem_246_3_W0_clk;
  wire [7:0] mem_246_3_W0_data;
  wire  mem_246_3_W0_en;
  wire  mem_246_3_W0_mask;
  wire [25:0] mem_246_4_R0_addr;
  wire  mem_246_4_R0_clk;
  wire [7:0] mem_246_4_R0_data;
  wire  mem_246_4_R0_en;
  wire [25:0] mem_246_4_W0_addr;
  wire  mem_246_4_W0_clk;
  wire [7:0] mem_246_4_W0_data;
  wire  mem_246_4_W0_en;
  wire  mem_246_4_W0_mask;
  wire [25:0] mem_246_5_R0_addr;
  wire  mem_246_5_R0_clk;
  wire [7:0] mem_246_5_R0_data;
  wire  mem_246_5_R0_en;
  wire [25:0] mem_246_5_W0_addr;
  wire  mem_246_5_W0_clk;
  wire [7:0] mem_246_5_W0_data;
  wire  mem_246_5_W0_en;
  wire  mem_246_5_W0_mask;
  wire [25:0] mem_246_6_R0_addr;
  wire  mem_246_6_R0_clk;
  wire [7:0] mem_246_6_R0_data;
  wire  mem_246_6_R0_en;
  wire [25:0] mem_246_6_W0_addr;
  wire  mem_246_6_W0_clk;
  wire [7:0] mem_246_6_W0_data;
  wire  mem_246_6_W0_en;
  wire  mem_246_6_W0_mask;
  wire [25:0] mem_246_7_R0_addr;
  wire  mem_246_7_R0_clk;
  wire [7:0] mem_246_7_R0_data;
  wire  mem_246_7_R0_en;
  wire [25:0] mem_246_7_W0_addr;
  wire  mem_246_7_W0_clk;
  wire [7:0] mem_246_7_W0_data;
  wire  mem_246_7_W0_en;
  wire  mem_246_7_W0_mask;
  wire [25:0] mem_247_0_R0_addr;
  wire  mem_247_0_R0_clk;
  wire [7:0] mem_247_0_R0_data;
  wire  mem_247_0_R0_en;
  wire [25:0] mem_247_0_W0_addr;
  wire  mem_247_0_W0_clk;
  wire [7:0] mem_247_0_W0_data;
  wire  mem_247_0_W0_en;
  wire  mem_247_0_W0_mask;
  wire [25:0] mem_247_1_R0_addr;
  wire  mem_247_1_R0_clk;
  wire [7:0] mem_247_1_R0_data;
  wire  mem_247_1_R0_en;
  wire [25:0] mem_247_1_W0_addr;
  wire  mem_247_1_W0_clk;
  wire [7:0] mem_247_1_W0_data;
  wire  mem_247_1_W0_en;
  wire  mem_247_1_W0_mask;
  wire [25:0] mem_247_2_R0_addr;
  wire  mem_247_2_R0_clk;
  wire [7:0] mem_247_2_R0_data;
  wire  mem_247_2_R0_en;
  wire [25:0] mem_247_2_W0_addr;
  wire  mem_247_2_W0_clk;
  wire [7:0] mem_247_2_W0_data;
  wire  mem_247_2_W0_en;
  wire  mem_247_2_W0_mask;
  wire [25:0] mem_247_3_R0_addr;
  wire  mem_247_3_R0_clk;
  wire [7:0] mem_247_3_R0_data;
  wire  mem_247_3_R0_en;
  wire [25:0] mem_247_3_W0_addr;
  wire  mem_247_3_W0_clk;
  wire [7:0] mem_247_3_W0_data;
  wire  mem_247_3_W0_en;
  wire  mem_247_3_W0_mask;
  wire [25:0] mem_247_4_R0_addr;
  wire  mem_247_4_R0_clk;
  wire [7:0] mem_247_4_R0_data;
  wire  mem_247_4_R0_en;
  wire [25:0] mem_247_4_W0_addr;
  wire  mem_247_4_W0_clk;
  wire [7:0] mem_247_4_W0_data;
  wire  mem_247_4_W0_en;
  wire  mem_247_4_W0_mask;
  wire [25:0] mem_247_5_R0_addr;
  wire  mem_247_5_R0_clk;
  wire [7:0] mem_247_5_R0_data;
  wire  mem_247_5_R0_en;
  wire [25:0] mem_247_5_W0_addr;
  wire  mem_247_5_W0_clk;
  wire [7:0] mem_247_5_W0_data;
  wire  mem_247_5_W0_en;
  wire  mem_247_5_W0_mask;
  wire [25:0] mem_247_6_R0_addr;
  wire  mem_247_6_R0_clk;
  wire [7:0] mem_247_6_R0_data;
  wire  mem_247_6_R0_en;
  wire [25:0] mem_247_6_W0_addr;
  wire  mem_247_6_W0_clk;
  wire [7:0] mem_247_6_W0_data;
  wire  mem_247_6_W0_en;
  wire  mem_247_6_W0_mask;
  wire [25:0] mem_247_7_R0_addr;
  wire  mem_247_7_R0_clk;
  wire [7:0] mem_247_7_R0_data;
  wire  mem_247_7_R0_en;
  wire [25:0] mem_247_7_W0_addr;
  wire  mem_247_7_W0_clk;
  wire [7:0] mem_247_7_W0_data;
  wire  mem_247_7_W0_en;
  wire  mem_247_7_W0_mask;
  wire [25:0] mem_248_0_R0_addr;
  wire  mem_248_0_R0_clk;
  wire [7:0] mem_248_0_R0_data;
  wire  mem_248_0_R0_en;
  wire [25:0] mem_248_0_W0_addr;
  wire  mem_248_0_W0_clk;
  wire [7:0] mem_248_0_W0_data;
  wire  mem_248_0_W0_en;
  wire  mem_248_0_W0_mask;
  wire [25:0] mem_248_1_R0_addr;
  wire  mem_248_1_R0_clk;
  wire [7:0] mem_248_1_R0_data;
  wire  mem_248_1_R0_en;
  wire [25:0] mem_248_1_W0_addr;
  wire  mem_248_1_W0_clk;
  wire [7:0] mem_248_1_W0_data;
  wire  mem_248_1_W0_en;
  wire  mem_248_1_W0_mask;
  wire [25:0] mem_248_2_R0_addr;
  wire  mem_248_2_R0_clk;
  wire [7:0] mem_248_2_R0_data;
  wire  mem_248_2_R0_en;
  wire [25:0] mem_248_2_W0_addr;
  wire  mem_248_2_W0_clk;
  wire [7:0] mem_248_2_W0_data;
  wire  mem_248_2_W0_en;
  wire  mem_248_2_W0_mask;
  wire [25:0] mem_248_3_R0_addr;
  wire  mem_248_3_R0_clk;
  wire [7:0] mem_248_3_R0_data;
  wire  mem_248_3_R0_en;
  wire [25:0] mem_248_3_W0_addr;
  wire  mem_248_3_W0_clk;
  wire [7:0] mem_248_3_W0_data;
  wire  mem_248_3_W0_en;
  wire  mem_248_3_W0_mask;
  wire [25:0] mem_248_4_R0_addr;
  wire  mem_248_4_R0_clk;
  wire [7:0] mem_248_4_R0_data;
  wire  mem_248_4_R0_en;
  wire [25:0] mem_248_4_W0_addr;
  wire  mem_248_4_W0_clk;
  wire [7:0] mem_248_4_W0_data;
  wire  mem_248_4_W0_en;
  wire  mem_248_4_W0_mask;
  wire [25:0] mem_248_5_R0_addr;
  wire  mem_248_5_R0_clk;
  wire [7:0] mem_248_5_R0_data;
  wire  mem_248_5_R0_en;
  wire [25:0] mem_248_5_W0_addr;
  wire  mem_248_5_W0_clk;
  wire [7:0] mem_248_5_W0_data;
  wire  mem_248_5_W0_en;
  wire  mem_248_5_W0_mask;
  wire [25:0] mem_248_6_R0_addr;
  wire  mem_248_6_R0_clk;
  wire [7:0] mem_248_6_R0_data;
  wire  mem_248_6_R0_en;
  wire [25:0] mem_248_6_W0_addr;
  wire  mem_248_6_W0_clk;
  wire [7:0] mem_248_6_W0_data;
  wire  mem_248_6_W0_en;
  wire  mem_248_6_W0_mask;
  wire [25:0] mem_248_7_R0_addr;
  wire  mem_248_7_R0_clk;
  wire [7:0] mem_248_7_R0_data;
  wire  mem_248_7_R0_en;
  wire [25:0] mem_248_7_W0_addr;
  wire  mem_248_7_W0_clk;
  wire [7:0] mem_248_7_W0_data;
  wire  mem_248_7_W0_en;
  wire  mem_248_7_W0_mask;
  wire [25:0] mem_249_0_R0_addr;
  wire  mem_249_0_R0_clk;
  wire [7:0] mem_249_0_R0_data;
  wire  mem_249_0_R0_en;
  wire [25:0] mem_249_0_W0_addr;
  wire  mem_249_0_W0_clk;
  wire [7:0] mem_249_0_W0_data;
  wire  mem_249_0_W0_en;
  wire  mem_249_0_W0_mask;
  wire [25:0] mem_249_1_R0_addr;
  wire  mem_249_1_R0_clk;
  wire [7:0] mem_249_1_R0_data;
  wire  mem_249_1_R0_en;
  wire [25:0] mem_249_1_W0_addr;
  wire  mem_249_1_W0_clk;
  wire [7:0] mem_249_1_W0_data;
  wire  mem_249_1_W0_en;
  wire  mem_249_1_W0_mask;
  wire [25:0] mem_249_2_R0_addr;
  wire  mem_249_2_R0_clk;
  wire [7:0] mem_249_2_R0_data;
  wire  mem_249_2_R0_en;
  wire [25:0] mem_249_2_W0_addr;
  wire  mem_249_2_W0_clk;
  wire [7:0] mem_249_2_W0_data;
  wire  mem_249_2_W0_en;
  wire  mem_249_2_W0_mask;
  wire [25:0] mem_249_3_R0_addr;
  wire  mem_249_3_R0_clk;
  wire [7:0] mem_249_3_R0_data;
  wire  mem_249_3_R0_en;
  wire [25:0] mem_249_3_W0_addr;
  wire  mem_249_3_W0_clk;
  wire [7:0] mem_249_3_W0_data;
  wire  mem_249_3_W0_en;
  wire  mem_249_3_W0_mask;
  wire [25:0] mem_249_4_R0_addr;
  wire  mem_249_4_R0_clk;
  wire [7:0] mem_249_4_R0_data;
  wire  mem_249_4_R0_en;
  wire [25:0] mem_249_4_W0_addr;
  wire  mem_249_4_W0_clk;
  wire [7:0] mem_249_4_W0_data;
  wire  mem_249_4_W0_en;
  wire  mem_249_4_W0_mask;
  wire [25:0] mem_249_5_R0_addr;
  wire  mem_249_5_R0_clk;
  wire [7:0] mem_249_5_R0_data;
  wire  mem_249_5_R0_en;
  wire [25:0] mem_249_5_W0_addr;
  wire  mem_249_5_W0_clk;
  wire [7:0] mem_249_5_W0_data;
  wire  mem_249_5_W0_en;
  wire  mem_249_5_W0_mask;
  wire [25:0] mem_249_6_R0_addr;
  wire  mem_249_6_R0_clk;
  wire [7:0] mem_249_6_R0_data;
  wire  mem_249_6_R0_en;
  wire [25:0] mem_249_6_W0_addr;
  wire  mem_249_6_W0_clk;
  wire [7:0] mem_249_6_W0_data;
  wire  mem_249_6_W0_en;
  wire  mem_249_6_W0_mask;
  wire [25:0] mem_249_7_R0_addr;
  wire  mem_249_7_R0_clk;
  wire [7:0] mem_249_7_R0_data;
  wire  mem_249_7_R0_en;
  wire [25:0] mem_249_7_W0_addr;
  wire  mem_249_7_W0_clk;
  wire [7:0] mem_249_7_W0_data;
  wire  mem_249_7_W0_en;
  wire  mem_249_7_W0_mask;
  wire [25:0] mem_250_0_R0_addr;
  wire  mem_250_0_R0_clk;
  wire [7:0] mem_250_0_R0_data;
  wire  mem_250_0_R0_en;
  wire [25:0] mem_250_0_W0_addr;
  wire  mem_250_0_W0_clk;
  wire [7:0] mem_250_0_W0_data;
  wire  mem_250_0_W0_en;
  wire  mem_250_0_W0_mask;
  wire [25:0] mem_250_1_R0_addr;
  wire  mem_250_1_R0_clk;
  wire [7:0] mem_250_1_R0_data;
  wire  mem_250_1_R0_en;
  wire [25:0] mem_250_1_W0_addr;
  wire  mem_250_1_W0_clk;
  wire [7:0] mem_250_1_W0_data;
  wire  mem_250_1_W0_en;
  wire  mem_250_1_W0_mask;
  wire [25:0] mem_250_2_R0_addr;
  wire  mem_250_2_R0_clk;
  wire [7:0] mem_250_2_R0_data;
  wire  mem_250_2_R0_en;
  wire [25:0] mem_250_2_W0_addr;
  wire  mem_250_2_W0_clk;
  wire [7:0] mem_250_2_W0_data;
  wire  mem_250_2_W0_en;
  wire  mem_250_2_W0_mask;
  wire [25:0] mem_250_3_R0_addr;
  wire  mem_250_3_R0_clk;
  wire [7:0] mem_250_3_R0_data;
  wire  mem_250_3_R0_en;
  wire [25:0] mem_250_3_W0_addr;
  wire  mem_250_3_W0_clk;
  wire [7:0] mem_250_3_W0_data;
  wire  mem_250_3_W0_en;
  wire  mem_250_3_W0_mask;
  wire [25:0] mem_250_4_R0_addr;
  wire  mem_250_4_R0_clk;
  wire [7:0] mem_250_4_R0_data;
  wire  mem_250_4_R0_en;
  wire [25:0] mem_250_4_W0_addr;
  wire  mem_250_4_W0_clk;
  wire [7:0] mem_250_4_W0_data;
  wire  mem_250_4_W0_en;
  wire  mem_250_4_W0_mask;
  wire [25:0] mem_250_5_R0_addr;
  wire  mem_250_5_R0_clk;
  wire [7:0] mem_250_5_R0_data;
  wire  mem_250_5_R0_en;
  wire [25:0] mem_250_5_W0_addr;
  wire  mem_250_5_W0_clk;
  wire [7:0] mem_250_5_W0_data;
  wire  mem_250_5_W0_en;
  wire  mem_250_5_W0_mask;
  wire [25:0] mem_250_6_R0_addr;
  wire  mem_250_6_R0_clk;
  wire [7:0] mem_250_6_R0_data;
  wire  mem_250_6_R0_en;
  wire [25:0] mem_250_6_W0_addr;
  wire  mem_250_6_W0_clk;
  wire [7:0] mem_250_6_W0_data;
  wire  mem_250_6_W0_en;
  wire  mem_250_6_W0_mask;
  wire [25:0] mem_250_7_R0_addr;
  wire  mem_250_7_R0_clk;
  wire [7:0] mem_250_7_R0_data;
  wire  mem_250_7_R0_en;
  wire [25:0] mem_250_7_W0_addr;
  wire  mem_250_7_W0_clk;
  wire [7:0] mem_250_7_W0_data;
  wire  mem_250_7_W0_en;
  wire  mem_250_7_W0_mask;
  wire [25:0] mem_251_0_R0_addr;
  wire  mem_251_0_R0_clk;
  wire [7:0] mem_251_0_R0_data;
  wire  mem_251_0_R0_en;
  wire [25:0] mem_251_0_W0_addr;
  wire  mem_251_0_W0_clk;
  wire [7:0] mem_251_0_W0_data;
  wire  mem_251_0_W0_en;
  wire  mem_251_0_W0_mask;
  wire [25:0] mem_251_1_R0_addr;
  wire  mem_251_1_R0_clk;
  wire [7:0] mem_251_1_R0_data;
  wire  mem_251_1_R0_en;
  wire [25:0] mem_251_1_W0_addr;
  wire  mem_251_1_W0_clk;
  wire [7:0] mem_251_1_W0_data;
  wire  mem_251_1_W0_en;
  wire  mem_251_1_W0_mask;
  wire [25:0] mem_251_2_R0_addr;
  wire  mem_251_2_R0_clk;
  wire [7:0] mem_251_2_R0_data;
  wire  mem_251_2_R0_en;
  wire [25:0] mem_251_2_W0_addr;
  wire  mem_251_2_W0_clk;
  wire [7:0] mem_251_2_W0_data;
  wire  mem_251_2_W0_en;
  wire  mem_251_2_W0_mask;
  wire [25:0] mem_251_3_R0_addr;
  wire  mem_251_3_R0_clk;
  wire [7:0] mem_251_3_R0_data;
  wire  mem_251_3_R0_en;
  wire [25:0] mem_251_3_W0_addr;
  wire  mem_251_3_W0_clk;
  wire [7:0] mem_251_3_W0_data;
  wire  mem_251_3_W0_en;
  wire  mem_251_3_W0_mask;
  wire [25:0] mem_251_4_R0_addr;
  wire  mem_251_4_R0_clk;
  wire [7:0] mem_251_4_R0_data;
  wire  mem_251_4_R0_en;
  wire [25:0] mem_251_4_W0_addr;
  wire  mem_251_4_W0_clk;
  wire [7:0] mem_251_4_W0_data;
  wire  mem_251_4_W0_en;
  wire  mem_251_4_W0_mask;
  wire [25:0] mem_251_5_R0_addr;
  wire  mem_251_5_R0_clk;
  wire [7:0] mem_251_5_R0_data;
  wire  mem_251_5_R0_en;
  wire [25:0] mem_251_5_W0_addr;
  wire  mem_251_5_W0_clk;
  wire [7:0] mem_251_5_W0_data;
  wire  mem_251_5_W0_en;
  wire  mem_251_5_W0_mask;
  wire [25:0] mem_251_6_R0_addr;
  wire  mem_251_6_R0_clk;
  wire [7:0] mem_251_6_R0_data;
  wire  mem_251_6_R0_en;
  wire [25:0] mem_251_6_W0_addr;
  wire  mem_251_6_W0_clk;
  wire [7:0] mem_251_6_W0_data;
  wire  mem_251_6_W0_en;
  wire  mem_251_6_W0_mask;
  wire [25:0] mem_251_7_R0_addr;
  wire  mem_251_7_R0_clk;
  wire [7:0] mem_251_7_R0_data;
  wire  mem_251_7_R0_en;
  wire [25:0] mem_251_7_W0_addr;
  wire  mem_251_7_W0_clk;
  wire [7:0] mem_251_7_W0_data;
  wire  mem_251_7_W0_en;
  wire  mem_251_7_W0_mask;
  wire [25:0] mem_252_0_R0_addr;
  wire  mem_252_0_R0_clk;
  wire [7:0] mem_252_0_R0_data;
  wire  mem_252_0_R0_en;
  wire [25:0] mem_252_0_W0_addr;
  wire  mem_252_0_W0_clk;
  wire [7:0] mem_252_0_W0_data;
  wire  mem_252_0_W0_en;
  wire  mem_252_0_W0_mask;
  wire [25:0] mem_252_1_R0_addr;
  wire  mem_252_1_R0_clk;
  wire [7:0] mem_252_1_R0_data;
  wire  mem_252_1_R0_en;
  wire [25:0] mem_252_1_W0_addr;
  wire  mem_252_1_W0_clk;
  wire [7:0] mem_252_1_W0_data;
  wire  mem_252_1_W0_en;
  wire  mem_252_1_W0_mask;
  wire [25:0] mem_252_2_R0_addr;
  wire  mem_252_2_R0_clk;
  wire [7:0] mem_252_2_R0_data;
  wire  mem_252_2_R0_en;
  wire [25:0] mem_252_2_W0_addr;
  wire  mem_252_2_W0_clk;
  wire [7:0] mem_252_2_W0_data;
  wire  mem_252_2_W0_en;
  wire  mem_252_2_W0_mask;
  wire [25:0] mem_252_3_R0_addr;
  wire  mem_252_3_R0_clk;
  wire [7:0] mem_252_3_R0_data;
  wire  mem_252_3_R0_en;
  wire [25:0] mem_252_3_W0_addr;
  wire  mem_252_3_W0_clk;
  wire [7:0] mem_252_3_W0_data;
  wire  mem_252_3_W0_en;
  wire  mem_252_3_W0_mask;
  wire [25:0] mem_252_4_R0_addr;
  wire  mem_252_4_R0_clk;
  wire [7:0] mem_252_4_R0_data;
  wire  mem_252_4_R0_en;
  wire [25:0] mem_252_4_W0_addr;
  wire  mem_252_4_W0_clk;
  wire [7:0] mem_252_4_W0_data;
  wire  mem_252_4_W0_en;
  wire  mem_252_4_W0_mask;
  wire [25:0] mem_252_5_R0_addr;
  wire  mem_252_5_R0_clk;
  wire [7:0] mem_252_5_R0_data;
  wire  mem_252_5_R0_en;
  wire [25:0] mem_252_5_W0_addr;
  wire  mem_252_5_W0_clk;
  wire [7:0] mem_252_5_W0_data;
  wire  mem_252_5_W0_en;
  wire  mem_252_5_W0_mask;
  wire [25:0] mem_252_6_R0_addr;
  wire  mem_252_6_R0_clk;
  wire [7:0] mem_252_6_R0_data;
  wire  mem_252_6_R0_en;
  wire [25:0] mem_252_6_W0_addr;
  wire  mem_252_6_W0_clk;
  wire [7:0] mem_252_6_W0_data;
  wire  mem_252_6_W0_en;
  wire  mem_252_6_W0_mask;
  wire [25:0] mem_252_7_R0_addr;
  wire  mem_252_7_R0_clk;
  wire [7:0] mem_252_7_R0_data;
  wire  mem_252_7_R0_en;
  wire [25:0] mem_252_7_W0_addr;
  wire  mem_252_7_W0_clk;
  wire [7:0] mem_252_7_W0_data;
  wire  mem_252_7_W0_en;
  wire  mem_252_7_W0_mask;
  wire [25:0] mem_253_0_R0_addr;
  wire  mem_253_0_R0_clk;
  wire [7:0] mem_253_0_R0_data;
  wire  mem_253_0_R0_en;
  wire [25:0] mem_253_0_W0_addr;
  wire  mem_253_0_W0_clk;
  wire [7:0] mem_253_0_W0_data;
  wire  mem_253_0_W0_en;
  wire  mem_253_0_W0_mask;
  wire [25:0] mem_253_1_R0_addr;
  wire  mem_253_1_R0_clk;
  wire [7:0] mem_253_1_R0_data;
  wire  mem_253_1_R0_en;
  wire [25:0] mem_253_1_W0_addr;
  wire  mem_253_1_W0_clk;
  wire [7:0] mem_253_1_W0_data;
  wire  mem_253_1_W0_en;
  wire  mem_253_1_W0_mask;
  wire [25:0] mem_253_2_R0_addr;
  wire  mem_253_2_R0_clk;
  wire [7:0] mem_253_2_R0_data;
  wire  mem_253_2_R0_en;
  wire [25:0] mem_253_2_W0_addr;
  wire  mem_253_2_W0_clk;
  wire [7:0] mem_253_2_W0_data;
  wire  mem_253_2_W0_en;
  wire  mem_253_2_W0_mask;
  wire [25:0] mem_253_3_R0_addr;
  wire  mem_253_3_R0_clk;
  wire [7:0] mem_253_3_R0_data;
  wire  mem_253_3_R0_en;
  wire [25:0] mem_253_3_W0_addr;
  wire  mem_253_3_W0_clk;
  wire [7:0] mem_253_3_W0_data;
  wire  mem_253_3_W0_en;
  wire  mem_253_3_W0_mask;
  wire [25:0] mem_253_4_R0_addr;
  wire  mem_253_4_R0_clk;
  wire [7:0] mem_253_4_R0_data;
  wire  mem_253_4_R0_en;
  wire [25:0] mem_253_4_W0_addr;
  wire  mem_253_4_W0_clk;
  wire [7:0] mem_253_4_W0_data;
  wire  mem_253_4_W0_en;
  wire  mem_253_4_W0_mask;
  wire [25:0] mem_253_5_R0_addr;
  wire  mem_253_5_R0_clk;
  wire [7:0] mem_253_5_R0_data;
  wire  mem_253_5_R0_en;
  wire [25:0] mem_253_5_W0_addr;
  wire  mem_253_5_W0_clk;
  wire [7:0] mem_253_5_W0_data;
  wire  mem_253_5_W0_en;
  wire  mem_253_5_W0_mask;
  wire [25:0] mem_253_6_R0_addr;
  wire  mem_253_6_R0_clk;
  wire [7:0] mem_253_6_R0_data;
  wire  mem_253_6_R0_en;
  wire [25:0] mem_253_6_W0_addr;
  wire  mem_253_6_W0_clk;
  wire [7:0] mem_253_6_W0_data;
  wire  mem_253_6_W0_en;
  wire  mem_253_6_W0_mask;
  wire [25:0] mem_253_7_R0_addr;
  wire  mem_253_7_R0_clk;
  wire [7:0] mem_253_7_R0_data;
  wire  mem_253_7_R0_en;
  wire [25:0] mem_253_7_W0_addr;
  wire  mem_253_7_W0_clk;
  wire [7:0] mem_253_7_W0_data;
  wire  mem_253_7_W0_en;
  wire  mem_253_7_W0_mask;
  wire [25:0] mem_254_0_R0_addr;
  wire  mem_254_0_R0_clk;
  wire [7:0] mem_254_0_R0_data;
  wire  mem_254_0_R0_en;
  wire [25:0] mem_254_0_W0_addr;
  wire  mem_254_0_W0_clk;
  wire [7:0] mem_254_0_W0_data;
  wire  mem_254_0_W0_en;
  wire  mem_254_0_W0_mask;
  wire [25:0] mem_254_1_R0_addr;
  wire  mem_254_1_R0_clk;
  wire [7:0] mem_254_1_R0_data;
  wire  mem_254_1_R0_en;
  wire [25:0] mem_254_1_W0_addr;
  wire  mem_254_1_W0_clk;
  wire [7:0] mem_254_1_W0_data;
  wire  mem_254_1_W0_en;
  wire  mem_254_1_W0_mask;
  wire [25:0] mem_254_2_R0_addr;
  wire  mem_254_2_R0_clk;
  wire [7:0] mem_254_2_R0_data;
  wire  mem_254_2_R0_en;
  wire [25:0] mem_254_2_W0_addr;
  wire  mem_254_2_W0_clk;
  wire [7:0] mem_254_2_W0_data;
  wire  mem_254_2_W0_en;
  wire  mem_254_2_W0_mask;
  wire [25:0] mem_254_3_R0_addr;
  wire  mem_254_3_R0_clk;
  wire [7:0] mem_254_3_R0_data;
  wire  mem_254_3_R0_en;
  wire [25:0] mem_254_3_W0_addr;
  wire  mem_254_3_W0_clk;
  wire [7:0] mem_254_3_W0_data;
  wire  mem_254_3_W0_en;
  wire  mem_254_3_W0_mask;
  wire [25:0] mem_254_4_R0_addr;
  wire  mem_254_4_R0_clk;
  wire [7:0] mem_254_4_R0_data;
  wire  mem_254_4_R0_en;
  wire [25:0] mem_254_4_W0_addr;
  wire  mem_254_4_W0_clk;
  wire [7:0] mem_254_4_W0_data;
  wire  mem_254_4_W0_en;
  wire  mem_254_4_W0_mask;
  wire [25:0] mem_254_5_R0_addr;
  wire  mem_254_5_R0_clk;
  wire [7:0] mem_254_5_R0_data;
  wire  mem_254_5_R0_en;
  wire [25:0] mem_254_5_W0_addr;
  wire  mem_254_5_W0_clk;
  wire [7:0] mem_254_5_W0_data;
  wire  mem_254_5_W0_en;
  wire  mem_254_5_W0_mask;
  wire [25:0] mem_254_6_R0_addr;
  wire  mem_254_6_R0_clk;
  wire [7:0] mem_254_6_R0_data;
  wire  mem_254_6_R0_en;
  wire [25:0] mem_254_6_W0_addr;
  wire  mem_254_6_W0_clk;
  wire [7:0] mem_254_6_W0_data;
  wire  mem_254_6_W0_en;
  wire  mem_254_6_W0_mask;
  wire [25:0] mem_254_7_R0_addr;
  wire  mem_254_7_R0_clk;
  wire [7:0] mem_254_7_R0_data;
  wire  mem_254_7_R0_en;
  wire [25:0] mem_254_7_W0_addr;
  wire  mem_254_7_W0_clk;
  wire [7:0] mem_254_7_W0_data;
  wire  mem_254_7_W0_en;
  wire  mem_254_7_W0_mask;
  wire [25:0] mem_255_0_R0_addr;
  wire  mem_255_0_R0_clk;
  wire [7:0] mem_255_0_R0_data;
  wire  mem_255_0_R0_en;
  wire [25:0] mem_255_0_W0_addr;
  wire  mem_255_0_W0_clk;
  wire [7:0] mem_255_0_W0_data;
  wire  mem_255_0_W0_en;
  wire  mem_255_0_W0_mask;
  wire [25:0] mem_255_1_R0_addr;
  wire  mem_255_1_R0_clk;
  wire [7:0] mem_255_1_R0_data;
  wire  mem_255_1_R0_en;
  wire [25:0] mem_255_1_W0_addr;
  wire  mem_255_1_W0_clk;
  wire [7:0] mem_255_1_W0_data;
  wire  mem_255_1_W0_en;
  wire  mem_255_1_W0_mask;
  wire [25:0] mem_255_2_R0_addr;
  wire  mem_255_2_R0_clk;
  wire [7:0] mem_255_2_R0_data;
  wire  mem_255_2_R0_en;
  wire [25:0] mem_255_2_W0_addr;
  wire  mem_255_2_W0_clk;
  wire [7:0] mem_255_2_W0_data;
  wire  mem_255_2_W0_en;
  wire  mem_255_2_W0_mask;
  wire [25:0] mem_255_3_R0_addr;
  wire  mem_255_3_R0_clk;
  wire [7:0] mem_255_3_R0_data;
  wire  mem_255_3_R0_en;
  wire [25:0] mem_255_3_W0_addr;
  wire  mem_255_3_W0_clk;
  wire [7:0] mem_255_3_W0_data;
  wire  mem_255_3_W0_en;
  wire  mem_255_3_W0_mask;
  wire [25:0] mem_255_4_R0_addr;
  wire  mem_255_4_R0_clk;
  wire [7:0] mem_255_4_R0_data;
  wire  mem_255_4_R0_en;
  wire [25:0] mem_255_4_W0_addr;
  wire  mem_255_4_W0_clk;
  wire [7:0] mem_255_4_W0_data;
  wire  mem_255_4_W0_en;
  wire  mem_255_4_W0_mask;
  wire [25:0] mem_255_5_R0_addr;
  wire  mem_255_5_R0_clk;
  wire [7:0] mem_255_5_R0_data;
  wire  mem_255_5_R0_en;
  wire [25:0] mem_255_5_W0_addr;
  wire  mem_255_5_W0_clk;
  wire [7:0] mem_255_5_W0_data;
  wire  mem_255_5_W0_en;
  wire  mem_255_5_W0_mask;
  wire [25:0] mem_255_6_R0_addr;
  wire  mem_255_6_R0_clk;
  wire [7:0] mem_255_6_R0_data;
  wire  mem_255_6_R0_en;
  wire [25:0] mem_255_6_W0_addr;
  wire  mem_255_6_W0_clk;
  wire [7:0] mem_255_6_W0_data;
  wire  mem_255_6_W0_en;
  wire  mem_255_6_W0_mask;
  wire [25:0] mem_255_7_R0_addr;
  wire  mem_255_7_R0_clk;
  wire [7:0] mem_255_7_R0_data;
  wire  mem_255_7_R0_en;
  wire [25:0] mem_255_7_W0_addr;
  wire  mem_255_7_W0_clk;
  wire [7:0] mem_255_7_W0_data;
  wire  mem_255_7_W0_en;
  wire  mem_255_7_W0_mask;
  wire [7:0] R0_addr_sel = R0_addr[33:26];
  reg [7:0] R0_addr_sel_reg;
  wire [7:0] W0_addr_sel = W0_addr[33:26];
  wire [7:0] R0_data_0_0 = mem_0_0_R0_data;
  wire [7:0] R0_data_0_1 = mem_0_1_R0_data;
  wire [7:0] R0_data_0_2 = mem_0_2_R0_data;
  wire [7:0] R0_data_0_3 = mem_0_3_R0_data;
  wire [7:0] R0_data_0_4 = mem_0_4_R0_data;
  wire [7:0] R0_data_0_5 = mem_0_5_R0_data;
  wire [7:0] R0_data_0_6 = mem_0_6_R0_data;
  wire [7:0] R0_data_0_7 = mem_0_7_R0_data;
  wire [63:0] R0_data_0 = {R0_data_0_7,R0_data_0_6,R0_data_0_5,R0_data_0_4,R0_data_0_3,R0_data_0_2,R0_data_0_1,
    R0_data_0_0};
  wire [7:0] R0_data_1_0 = mem_1_0_R0_data;
  wire [7:0] R0_data_1_1 = mem_1_1_R0_data;
  wire [7:0] R0_data_1_2 = mem_1_2_R0_data;
  wire [7:0] R0_data_1_3 = mem_1_3_R0_data;
  wire [7:0] R0_data_1_4 = mem_1_4_R0_data;
  wire [7:0] R0_data_1_5 = mem_1_5_R0_data;
  wire [7:0] R0_data_1_6 = mem_1_6_R0_data;
  wire [7:0] R0_data_1_7 = mem_1_7_R0_data;
  wire [63:0] R0_data_1 = {R0_data_1_7,R0_data_1_6,R0_data_1_5,R0_data_1_4,R0_data_1_3,R0_data_1_2,R0_data_1_1,
    R0_data_1_0};
  wire [7:0] R0_data_2_0 = mem_2_0_R0_data;
  wire [7:0] R0_data_2_1 = mem_2_1_R0_data;
  wire [7:0] R0_data_2_2 = mem_2_2_R0_data;
  wire [7:0] R0_data_2_3 = mem_2_3_R0_data;
  wire [7:0] R0_data_2_4 = mem_2_4_R0_data;
  wire [7:0] R0_data_2_5 = mem_2_5_R0_data;
  wire [7:0] R0_data_2_6 = mem_2_6_R0_data;
  wire [7:0] R0_data_2_7 = mem_2_7_R0_data;
  wire [63:0] R0_data_2 = {R0_data_2_7,R0_data_2_6,R0_data_2_5,R0_data_2_4,R0_data_2_3,R0_data_2_2,R0_data_2_1,
    R0_data_2_0};
  wire [7:0] R0_data_3_0 = mem_3_0_R0_data;
  wire [7:0] R0_data_3_1 = mem_3_1_R0_data;
  wire [7:0] R0_data_3_2 = mem_3_2_R0_data;
  wire [7:0] R0_data_3_3 = mem_3_3_R0_data;
  wire [7:0] R0_data_3_4 = mem_3_4_R0_data;
  wire [7:0] R0_data_3_5 = mem_3_5_R0_data;
  wire [7:0] R0_data_3_6 = mem_3_6_R0_data;
  wire [7:0] R0_data_3_7 = mem_3_7_R0_data;
  wire [63:0] R0_data_3 = {R0_data_3_7,R0_data_3_6,R0_data_3_5,R0_data_3_4,R0_data_3_3,R0_data_3_2,R0_data_3_1,
    R0_data_3_0};
  wire [7:0] R0_data_4_0 = mem_4_0_R0_data;
  wire [7:0] R0_data_4_1 = mem_4_1_R0_data;
  wire [7:0] R0_data_4_2 = mem_4_2_R0_data;
  wire [7:0] R0_data_4_3 = mem_4_3_R0_data;
  wire [7:0] R0_data_4_4 = mem_4_4_R0_data;
  wire [7:0] R0_data_4_5 = mem_4_5_R0_data;
  wire [7:0] R0_data_4_6 = mem_4_6_R0_data;
  wire [7:0] R0_data_4_7 = mem_4_7_R0_data;
  wire [63:0] R0_data_4 = {R0_data_4_7,R0_data_4_6,R0_data_4_5,R0_data_4_4,R0_data_4_3,R0_data_4_2,R0_data_4_1,
    R0_data_4_0};
  wire [7:0] R0_data_5_0 = mem_5_0_R0_data;
  wire [7:0] R0_data_5_1 = mem_5_1_R0_data;
  wire [7:0] R0_data_5_2 = mem_5_2_R0_data;
  wire [7:0] R0_data_5_3 = mem_5_3_R0_data;
  wire [7:0] R0_data_5_4 = mem_5_4_R0_data;
  wire [7:0] R0_data_5_5 = mem_5_5_R0_data;
  wire [7:0] R0_data_5_6 = mem_5_6_R0_data;
  wire [7:0] R0_data_5_7 = mem_5_7_R0_data;
  wire [63:0] R0_data_5 = {R0_data_5_7,R0_data_5_6,R0_data_5_5,R0_data_5_4,R0_data_5_3,R0_data_5_2,R0_data_5_1,
    R0_data_5_0};
  wire [7:0] R0_data_6_0 = mem_6_0_R0_data;
  wire [7:0] R0_data_6_1 = mem_6_1_R0_data;
  wire [7:0] R0_data_6_2 = mem_6_2_R0_data;
  wire [7:0] R0_data_6_3 = mem_6_3_R0_data;
  wire [7:0] R0_data_6_4 = mem_6_4_R0_data;
  wire [7:0] R0_data_6_5 = mem_6_5_R0_data;
  wire [7:0] R0_data_6_6 = mem_6_6_R0_data;
  wire [7:0] R0_data_6_7 = mem_6_7_R0_data;
  wire [63:0] R0_data_6 = {R0_data_6_7,R0_data_6_6,R0_data_6_5,R0_data_6_4,R0_data_6_3,R0_data_6_2,R0_data_6_1,
    R0_data_6_0};
  wire [7:0] R0_data_7_0 = mem_7_0_R0_data;
  wire [7:0] R0_data_7_1 = mem_7_1_R0_data;
  wire [7:0] R0_data_7_2 = mem_7_2_R0_data;
  wire [7:0] R0_data_7_3 = mem_7_3_R0_data;
  wire [7:0] R0_data_7_4 = mem_7_4_R0_data;
  wire [7:0] R0_data_7_5 = mem_7_5_R0_data;
  wire [7:0] R0_data_7_6 = mem_7_6_R0_data;
  wire [7:0] R0_data_7_7 = mem_7_7_R0_data;
  wire [63:0] R0_data_7 = {R0_data_7_7,R0_data_7_6,R0_data_7_5,R0_data_7_4,R0_data_7_3,R0_data_7_2,R0_data_7_1,
    R0_data_7_0};
  wire [7:0] R0_data_8_0 = mem_8_0_R0_data;
  wire [7:0] R0_data_8_1 = mem_8_1_R0_data;
  wire [7:0] R0_data_8_2 = mem_8_2_R0_data;
  wire [7:0] R0_data_8_3 = mem_8_3_R0_data;
  wire [7:0] R0_data_8_4 = mem_8_4_R0_data;
  wire [7:0] R0_data_8_5 = mem_8_5_R0_data;
  wire [7:0] R0_data_8_6 = mem_8_6_R0_data;
  wire [7:0] R0_data_8_7 = mem_8_7_R0_data;
  wire [63:0] R0_data_8 = {R0_data_8_7,R0_data_8_6,R0_data_8_5,R0_data_8_4,R0_data_8_3,R0_data_8_2,R0_data_8_1,
    R0_data_8_0};
  wire [7:0] R0_data_9_0 = mem_9_0_R0_data;
  wire [7:0] R0_data_9_1 = mem_9_1_R0_data;
  wire [7:0] R0_data_9_2 = mem_9_2_R0_data;
  wire [7:0] R0_data_9_3 = mem_9_3_R0_data;
  wire [7:0] R0_data_9_4 = mem_9_4_R0_data;
  wire [7:0] R0_data_9_5 = mem_9_5_R0_data;
  wire [7:0] R0_data_9_6 = mem_9_6_R0_data;
  wire [7:0] R0_data_9_7 = mem_9_7_R0_data;
  wire [63:0] R0_data_9 = {R0_data_9_7,R0_data_9_6,R0_data_9_5,R0_data_9_4,R0_data_9_3,R0_data_9_2,R0_data_9_1,
    R0_data_9_0};
  wire [7:0] R0_data_10_0 = mem_10_0_R0_data;
  wire [7:0] R0_data_10_1 = mem_10_1_R0_data;
  wire [7:0] R0_data_10_2 = mem_10_2_R0_data;
  wire [7:0] R0_data_10_3 = mem_10_3_R0_data;
  wire [7:0] R0_data_10_4 = mem_10_4_R0_data;
  wire [7:0] R0_data_10_5 = mem_10_5_R0_data;
  wire [7:0] R0_data_10_6 = mem_10_6_R0_data;
  wire [7:0] R0_data_10_7 = mem_10_7_R0_data;
  wire [63:0] R0_data_10 = {R0_data_10_7,R0_data_10_6,R0_data_10_5,R0_data_10_4,R0_data_10_3,R0_data_10_2,R0_data_10_1,
    R0_data_10_0};
  wire [7:0] R0_data_11_0 = mem_11_0_R0_data;
  wire [7:0] R0_data_11_1 = mem_11_1_R0_data;
  wire [7:0] R0_data_11_2 = mem_11_2_R0_data;
  wire [7:0] R0_data_11_3 = mem_11_3_R0_data;
  wire [7:0] R0_data_11_4 = mem_11_4_R0_data;
  wire [7:0] R0_data_11_5 = mem_11_5_R0_data;
  wire [7:0] R0_data_11_6 = mem_11_6_R0_data;
  wire [7:0] R0_data_11_7 = mem_11_7_R0_data;
  wire [63:0] R0_data_11 = {R0_data_11_7,R0_data_11_6,R0_data_11_5,R0_data_11_4,R0_data_11_3,R0_data_11_2,R0_data_11_1,
    R0_data_11_0};
  wire [7:0] R0_data_12_0 = mem_12_0_R0_data;
  wire [7:0] R0_data_12_1 = mem_12_1_R0_data;
  wire [7:0] R0_data_12_2 = mem_12_2_R0_data;
  wire [7:0] R0_data_12_3 = mem_12_3_R0_data;
  wire [7:0] R0_data_12_4 = mem_12_4_R0_data;
  wire [7:0] R0_data_12_5 = mem_12_5_R0_data;
  wire [7:0] R0_data_12_6 = mem_12_6_R0_data;
  wire [7:0] R0_data_12_7 = mem_12_7_R0_data;
  wire [63:0] R0_data_12 = {R0_data_12_7,R0_data_12_6,R0_data_12_5,R0_data_12_4,R0_data_12_3,R0_data_12_2,R0_data_12_1,
    R0_data_12_0};
  wire [7:0] R0_data_13_0 = mem_13_0_R0_data;
  wire [7:0] R0_data_13_1 = mem_13_1_R0_data;
  wire [7:0] R0_data_13_2 = mem_13_2_R0_data;
  wire [7:0] R0_data_13_3 = mem_13_3_R0_data;
  wire [7:0] R0_data_13_4 = mem_13_4_R0_data;
  wire [7:0] R0_data_13_5 = mem_13_5_R0_data;
  wire [7:0] R0_data_13_6 = mem_13_6_R0_data;
  wire [7:0] R0_data_13_7 = mem_13_7_R0_data;
  wire [63:0] R0_data_13 = {R0_data_13_7,R0_data_13_6,R0_data_13_5,R0_data_13_4,R0_data_13_3,R0_data_13_2,R0_data_13_1,
    R0_data_13_0};
  wire [7:0] R0_data_14_0 = mem_14_0_R0_data;
  wire [7:0] R0_data_14_1 = mem_14_1_R0_data;
  wire [7:0] R0_data_14_2 = mem_14_2_R0_data;
  wire [7:0] R0_data_14_3 = mem_14_3_R0_data;
  wire [7:0] R0_data_14_4 = mem_14_4_R0_data;
  wire [7:0] R0_data_14_5 = mem_14_5_R0_data;
  wire [7:0] R0_data_14_6 = mem_14_6_R0_data;
  wire [7:0] R0_data_14_7 = mem_14_7_R0_data;
  wire [63:0] R0_data_14 = {R0_data_14_7,R0_data_14_6,R0_data_14_5,R0_data_14_4,R0_data_14_3,R0_data_14_2,R0_data_14_1,
    R0_data_14_0};
  wire [7:0] R0_data_15_0 = mem_15_0_R0_data;
  wire [7:0] R0_data_15_1 = mem_15_1_R0_data;
  wire [7:0] R0_data_15_2 = mem_15_2_R0_data;
  wire [7:0] R0_data_15_3 = mem_15_3_R0_data;
  wire [7:0] R0_data_15_4 = mem_15_4_R0_data;
  wire [7:0] R0_data_15_5 = mem_15_5_R0_data;
  wire [7:0] R0_data_15_6 = mem_15_6_R0_data;
  wire [7:0] R0_data_15_7 = mem_15_7_R0_data;
  wire [63:0] R0_data_15 = {R0_data_15_7,R0_data_15_6,R0_data_15_5,R0_data_15_4,R0_data_15_3,R0_data_15_2,R0_data_15_1,
    R0_data_15_0};
  wire [7:0] R0_data_16_0 = mem_16_0_R0_data;
  wire [7:0] R0_data_16_1 = mem_16_1_R0_data;
  wire [7:0] R0_data_16_2 = mem_16_2_R0_data;
  wire [7:0] R0_data_16_3 = mem_16_3_R0_data;
  wire [7:0] R0_data_16_4 = mem_16_4_R0_data;
  wire [7:0] R0_data_16_5 = mem_16_5_R0_data;
  wire [7:0] R0_data_16_6 = mem_16_6_R0_data;
  wire [7:0] R0_data_16_7 = mem_16_7_R0_data;
  wire [63:0] R0_data_16 = {R0_data_16_7,R0_data_16_6,R0_data_16_5,R0_data_16_4,R0_data_16_3,R0_data_16_2,R0_data_16_1,
    R0_data_16_0};
  wire [7:0] R0_data_17_0 = mem_17_0_R0_data;
  wire [7:0] R0_data_17_1 = mem_17_1_R0_data;
  wire [7:0] R0_data_17_2 = mem_17_2_R0_data;
  wire [7:0] R0_data_17_3 = mem_17_3_R0_data;
  wire [7:0] R0_data_17_4 = mem_17_4_R0_data;
  wire [7:0] R0_data_17_5 = mem_17_5_R0_data;
  wire [7:0] R0_data_17_6 = mem_17_6_R0_data;
  wire [7:0] R0_data_17_7 = mem_17_7_R0_data;
  wire [63:0] R0_data_17 = {R0_data_17_7,R0_data_17_6,R0_data_17_5,R0_data_17_4,R0_data_17_3,R0_data_17_2,R0_data_17_1,
    R0_data_17_0};
  wire [7:0] R0_data_18_0 = mem_18_0_R0_data;
  wire [7:0] R0_data_18_1 = mem_18_1_R0_data;
  wire [7:0] R0_data_18_2 = mem_18_2_R0_data;
  wire [7:0] R0_data_18_3 = mem_18_3_R0_data;
  wire [7:0] R0_data_18_4 = mem_18_4_R0_data;
  wire [7:0] R0_data_18_5 = mem_18_5_R0_data;
  wire [7:0] R0_data_18_6 = mem_18_6_R0_data;
  wire [7:0] R0_data_18_7 = mem_18_7_R0_data;
  wire [63:0] R0_data_18 = {R0_data_18_7,R0_data_18_6,R0_data_18_5,R0_data_18_4,R0_data_18_3,R0_data_18_2,R0_data_18_1,
    R0_data_18_0};
  wire [7:0] R0_data_19_0 = mem_19_0_R0_data;
  wire [7:0] R0_data_19_1 = mem_19_1_R0_data;
  wire [7:0] R0_data_19_2 = mem_19_2_R0_data;
  wire [7:0] R0_data_19_3 = mem_19_3_R0_data;
  wire [7:0] R0_data_19_4 = mem_19_4_R0_data;
  wire [7:0] R0_data_19_5 = mem_19_5_R0_data;
  wire [7:0] R0_data_19_6 = mem_19_6_R0_data;
  wire [7:0] R0_data_19_7 = mem_19_7_R0_data;
  wire [63:0] R0_data_19 = {R0_data_19_7,R0_data_19_6,R0_data_19_5,R0_data_19_4,R0_data_19_3,R0_data_19_2,R0_data_19_1,
    R0_data_19_0};
  wire [7:0] R0_data_20_0 = mem_20_0_R0_data;
  wire [7:0] R0_data_20_1 = mem_20_1_R0_data;
  wire [7:0] R0_data_20_2 = mem_20_2_R0_data;
  wire [7:0] R0_data_20_3 = mem_20_3_R0_data;
  wire [7:0] R0_data_20_4 = mem_20_4_R0_data;
  wire [7:0] R0_data_20_5 = mem_20_5_R0_data;
  wire [7:0] R0_data_20_6 = mem_20_6_R0_data;
  wire [7:0] R0_data_20_7 = mem_20_7_R0_data;
  wire [63:0] R0_data_20 = {R0_data_20_7,R0_data_20_6,R0_data_20_5,R0_data_20_4,R0_data_20_3,R0_data_20_2,R0_data_20_1,
    R0_data_20_0};
  wire [7:0] R0_data_21_0 = mem_21_0_R0_data;
  wire [7:0] R0_data_21_1 = mem_21_1_R0_data;
  wire [7:0] R0_data_21_2 = mem_21_2_R0_data;
  wire [7:0] R0_data_21_3 = mem_21_3_R0_data;
  wire [7:0] R0_data_21_4 = mem_21_4_R0_data;
  wire [7:0] R0_data_21_5 = mem_21_5_R0_data;
  wire [7:0] R0_data_21_6 = mem_21_6_R0_data;
  wire [7:0] R0_data_21_7 = mem_21_7_R0_data;
  wire [63:0] R0_data_21 = {R0_data_21_7,R0_data_21_6,R0_data_21_5,R0_data_21_4,R0_data_21_3,R0_data_21_2,R0_data_21_1,
    R0_data_21_0};
  wire [7:0] R0_data_22_0 = mem_22_0_R0_data;
  wire [7:0] R0_data_22_1 = mem_22_1_R0_data;
  wire [7:0] R0_data_22_2 = mem_22_2_R0_data;
  wire [7:0] R0_data_22_3 = mem_22_3_R0_data;
  wire [7:0] R0_data_22_4 = mem_22_4_R0_data;
  wire [7:0] R0_data_22_5 = mem_22_5_R0_data;
  wire [7:0] R0_data_22_6 = mem_22_6_R0_data;
  wire [7:0] R0_data_22_7 = mem_22_7_R0_data;
  wire [63:0] R0_data_22 = {R0_data_22_7,R0_data_22_6,R0_data_22_5,R0_data_22_4,R0_data_22_3,R0_data_22_2,R0_data_22_1,
    R0_data_22_0};
  wire [7:0] R0_data_23_0 = mem_23_0_R0_data;
  wire [7:0] R0_data_23_1 = mem_23_1_R0_data;
  wire [7:0] R0_data_23_2 = mem_23_2_R0_data;
  wire [7:0] R0_data_23_3 = mem_23_3_R0_data;
  wire [7:0] R0_data_23_4 = mem_23_4_R0_data;
  wire [7:0] R0_data_23_5 = mem_23_5_R0_data;
  wire [7:0] R0_data_23_6 = mem_23_6_R0_data;
  wire [7:0] R0_data_23_7 = mem_23_7_R0_data;
  wire [63:0] R0_data_23 = {R0_data_23_7,R0_data_23_6,R0_data_23_5,R0_data_23_4,R0_data_23_3,R0_data_23_2,R0_data_23_1,
    R0_data_23_0};
  wire [7:0] R0_data_24_0 = mem_24_0_R0_data;
  wire [7:0] R0_data_24_1 = mem_24_1_R0_data;
  wire [7:0] R0_data_24_2 = mem_24_2_R0_data;
  wire [7:0] R0_data_24_3 = mem_24_3_R0_data;
  wire [7:0] R0_data_24_4 = mem_24_4_R0_data;
  wire [7:0] R0_data_24_5 = mem_24_5_R0_data;
  wire [7:0] R0_data_24_6 = mem_24_6_R0_data;
  wire [7:0] R0_data_24_7 = mem_24_7_R0_data;
  wire [63:0] R0_data_24 = {R0_data_24_7,R0_data_24_6,R0_data_24_5,R0_data_24_4,R0_data_24_3,R0_data_24_2,R0_data_24_1,
    R0_data_24_0};
  wire [7:0] R0_data_25_0 = mem_25_0_R0_data;
  wire [7:0] R0_data_25_1 = mem_25_1_R0_data;
  wire [7:0] R0_data_25_2 = mem_25_2_R0_data;
  wire [7:0] R0_data_25_3 = mem_25_3_R0_data;
  wire [7:0] R0_data_25_4 = mem_25_4_R0_data;
  wire [7:0] R0_data_25_5 = mem_25_5_R0_data;
  wire [7:0] R0_data_25_6 = mem_25_6_R0_data;
  wire [7:0] R0_data_25_7 = mem_25_7_R0_data;
  wire [63:0] R0_data_25 = {R0_data_25_7,R0_data_25_6,R0_data_25_5,R0_data_25_4,R0_data_25_3,R0_data_25_2,R0_data_25_1,
    R0_data_25_0};
  wire [7:0] R0_data_26_0 = mem_26_0_R0_data;
  wire [7:0] R0_data_26_1 = mem_26_1_R0_data;
  wire [7:0] R0_data_26_2 = mem_26_2_R0_data;
  wire [7:0] R0_data_26_3 = mem_26_3_R0_data;
  wire [7:0] R0_data_26_4 = mem_26_4_R0_data;
  wire [7:0] R0_data_26_5 = mem_26_5_R0_data;
  wire [7:0] R0_data_26_6 = mem_26_6_R0_data;
  wire [7:0] R0_data_26_7 = mem_26_7_R0_data;
  wire [63:0] R0_data_26 = {R0_data_26_7,R0_data_26_6,R0_data_26_5,R0_data_26_4,R0_data_26_3,R0_data_26_2,R0_data_26_1,
    R0_data_26_0};
  wire [7:0] R0_data_27_0 = mem_27_0_R0_data;
  wire [7:0] R0_data_27_1 = mem_27_1_R0_data;
  wire [7:0] R0_data_27_2 = mem_27_2_R0_data;
  wire [7:0] R0_data_27_3 = mem_27_3_R0_data;
  wire [7:0] R0_data_27_4 = mem_27_4_R0_data;
  wire [7:0] R0_data_27_5 = mem_27_5_R0_data;
  wire [7:0] R0_data_27_6 = mem_27_6_R0_data;
  wire [7:0] R0_data_27_7 = mem_27_7_R0_data;
  wire [63:0] R0_data_27 = {R0_data_27_7,R0_data_27_6,R0_data_27_5,R0_data_27_4,R0_data_27_3,R0_data_27_2,R0_data_27_1,
    R0_data_27_0};
  wire [7:0] R0_data_28_0 = mem_28_0_R0_data;
  wire [7:0] R0_data_28_1 = mem_28_1_R0_data;
  wire [7:0] R0_data_28_2 = mem_28_2_R0_data;
  wire [7:0] R0_data_28_3 = mem_28_3_R0_data;
  wire [7:0] R0_data_28_4 = mem_28_4_R0_data;
  wire [7:0] R0_data_28_5 = mem_28_5_R0_data;
  wire [7:0] R0_data_28_6 = mem_28_6_R0_data;
  wire [7:0] R0_data_28_7 = mem_28_7_R0_data;
  wire [63:0] R0_data_28 = {R0_data_28_7,R0_data_28_6,R0_data_28_5,R0_data_28_4,R0_data_28_3,R0_data_28_2,R0_data_28_1,
    R0_data_28_0};
  wire [7:0] R0_data_29_0 = mem_29_0_R0_data;
  wire [7:0] R0_data_29_1 = mem_29_1_R0_data;
  wire [7:0] R0_data_29_2 = mem_29_2_R0_data;
  wire [7:0] R0_data_29_3 = mem_29_3_R0_data;
  wire [7:0] R0_data_29_4 = mem_29_4_R0_data;
  wire [7:0] R0_data_29_5 = mem_29_5_R0_data;
  wire [7:0] R0_data_29_6 = mem_29_6_R0_data;
  wire [7:0] R0_data_29_7 = mem_29_7_R0_data;
  wire [63:0] R0_data_29 = {R0_data_29_7,R0_data_29_6,R0_data_29_5,R0_data_29_4,R0_data_29_3,R0_data_29_2,R0_data_29_1,
    R0_data_29_0};
  wire [7:0] R0_data_30_0 = mem_30_0_R0_data;
  wire [7:0] R0_data_30_1 = mem_30_1_R0_data;
  wire [7:0] R0_data_30_2 = mem_30_2_R0_data;
  wire [7:0] R0_data_30_3 = mem_30_3_R0_data;
  wire [7:0] R0_data_30_4 = mem_30_4_R0_data;
  wire [7:0] R0_data_30_5 = mem_30_5_R0_data;
  wire [7:0] R0_data_30_6 = mem_30_6_R0_data;
  wire [7:0] R0_data_30_7 = mem_30_7_R0_data;
  wire [63:0] R0_data_30 = {R0_data_30_7,R0_data_30_6,R0_data_30_5,R0_data_30_4,R0_data_30_3,R0_data_30_2,R0_data_30_1,
    R0_data_30_0};
  wire [7:0] R0_data_31_0 = mem_31_0_R0_data;
  wire [7:0] R0_data_31_1 = mem_31_1_R0_data;
  wire [7:0] R0_data_31_2 = mem_31_2_R0_data;
  wire [7:0] R0_data_31_3 = mem_31_3_R0_data;
  wire [7:0] R0_data_31_4 = mem_31_4_R0_data;
  wire [7:0] R0_data_31_5 = mem_31_5_R0_data;
  wire [7:0] R0_data_31_6 = mem_31_6_R0_data;
  wire [7:0] R0_data_31_7 = mem_31_7_R0_data;
  wire [63:0] R0_data_31 = {R0_data_31_7,R0_data_31_6,R0_data_31_5,R0_data_31_4,R0_data_31_3,R0_data_31_2,R0_data_31_1,
    R0_data_31_0};
  wire [7:0] R0_data_32_0 = mem_32_0_R0_data;
  wire [7:0] R0_data_32_1 = mem_32_1_R0_data;
  wire [7:0] R0_data_32_2 = mem_32_2_R0_data;
  wire [7:0] R0_data_32_3 = mem_32_3_R0_data;
  wire [7:0] R0_data_32_4 = mem_32_4_R0_data;
  wire [7:0] R0_data_32_5 = mem_32_5_R0_data;
  wire [7:0] R0_data_32_6 = mem_32_6_R0_data;
  wire [7:0] R0_data_32_7 = mem_32_7_R0_data;
  wire [63:0] R0_data_32 = {R0_data_32_7,R0_data_32_6,R0_data_32_5,R0_data_32_4,R0_data_32_3,R0_data_32_2,R0_data_32_1,
    R0_data_32_0};
  wire [7:0] R0_data_33_0 = mem_33_0_R0_data;
  wire [7:0] R0_data_33_1 = mem_33_1_R0_data;
  wire [7:0] R0_data_33_2 = mem_33_2_R0_data;
  wire [7:0] R0_data_33_3 = mem_33_3_R0_data;
  wire [7:0] R0_data_33_4 = mem_33_4_R0_data;
  wire [7:0] R0_data_33_5 = mem_33_5_R0_data;
  wire [7:0] R0_data_33_6 = mem_33_6_R0_data;
  wire [7:0] R0_data_33_7 = mem_33_7_R0_data;
  wire [63:0] R0_data_33 = {R0_data_33_7,R0_data_33_6,R0_data_33_5,R0_data_33_4,R0_data_33_3,R0_data_33_2,R0_data_33_1,
    R0_data_33_0};
  wire [7:0] R0_data_34_0 = mem_34_0_R0_data;
  wire [7:0] R0_data_34_1 = mem_34_1_R0_data;
  wire [7:0] R0_data_34_2 = mem_34_2_R0_data;
  wire [7:0] R0_data_34_3 = mem_34_3_R0_data;
  wire [7:0] R0_data_34_4 = mem_34_4_R0_data;
  wire [7:0] R0_data_34_5 = mem_34_5_R0_data;
  wire [7:0] R0_data_34_6 = mem_34_6_R0_data;
  wire [7:0] R0_data_34_7 = mem_34_7_R0_data;
  wire [63:0] R0_data_34 = {R0_data_34_7,R0_data_34_6,R0_data_34_5,R0_data_34_4,R0_data_34_3,R0_data_34_2,R0_data_34_1,
    R0_data_34_0};
  wire [7:0] R0_data_35_0 = mem_35_0_R0_data;
  wire [7:0] R0_data_35_1 = mem_35_1_R0_data;
  wire [7:0] R0_data_35_2 = mem_35_2_R0_data;
  wire [7:0] R0_data_35_3 = mem_35_3_R0_data;
  wire [7:0] R0_data_35_4 = mem_35_4_R0_data;
  wire [7:0] R0_data_35_5 = mem_35_5_R0_data;
  wire [7:0] R0_data_35_6 = mem_35_6_R0_data;
  wire [7:0] R0_data_35_7 = mem_35_7_R0_data;
  wire [63:0] R0_data_35 = {R0_data_35_7,R0_data_35_6,R0_data_35_5,R0_data_35_4,R0_data_35_3,R0_data_35_2,R0_data_35_1,
    R0_data_35_0};
  wire [7:0] R0_data_36_0 = mem_36_0_R0_data;
  wire [7:0] R0_data_36_1 = mem_36_1_R0_data;
  wire [7:0] R0_data_36_2 = mem_36_2_R0_data;
  wire [7:0] R0_data_36_3 = mem_36_3_R0_data;
  wire [7:0] R0_data_36_4 = mem_36_4_R0_data;
  wire [7:0] R0_data_36_5 = mem_36_5_R0_data;
  wire [7:0] R0_data_36_6 = mem_36_6_R0_data;
  wire [7:0] R0_data_36_7 = mem_36_7_R0_data;
  wire [63:0] R0_data_36 = {R0_data_36_7,R0_data_36_6,R0_data_36_5,R0_data_36_4,R0_data_36_3,R0_data_36_2,R0_data_36_1,
    R0_data_36_0};
  wire [7:0] R0_data_37_0 = mem_37_0_R0_data;
  wire [7:0] R0_data_37_1 = mem_37_1_R0_data;
  wire [7:0] R0_data_37_2 = mem_37_2_R0_data;
  wire [7:0] R0_data_37_3 = mem_37_3_R0_data;
  wire [7:0] R0_data_37_4 = mem_37_4_R0_data;
  wire [7:0] R0_data_37_5 = mem_37_5_R0_data;
  wire [7:0] R0_data_37_6 = mem_37_6_R0_data;
  wire [7:0] R0_data_37_7 = mem_37_7_R0_data;
  wire [63:0] R0_data_37 = {R0_data_37_7,R0_data_37_6,R0_data_37_5,R0_data_37_4,R0_data_37_3,R0_data_37_2,R0_data_37_1,
    R0_data_37_0};
  wire [7:0] R0_data_38_0 = mem_38_0_R0_data;
  wire [7:0] R0_data_38_1 = mem_38_1_R0_data;
  wire [7:0] R0_data_38_2 = mem_38_2_R0_data;
  wire [7:0] R0_data_38_3 = mem_38_3_R0_data;
  wire [7:0] R0_data_38_4 = mem_38_4_R0_data;
  wire [7:0] R0_data_38_5 = mem_38_5_R0_data;
  wire [7:0] R0_data_38_6 = mem_38_6_R0_data;
  wire [7:0] R0_data_38_7 = mem_38_7_R0_data;
  wire [63:0] R0_data_38 = {R0_data_38_7,R0_data_38_6,R0_data_38_5,R0_data_38_4,R0_data_38_3,R0_data_38_2,R0_data_38_1,
    R0_data_38_0};
  wire [7:0] R0_data_39_0 = mem_39_0_R0_data;
  wire [7:0] R0_data_39_1 = mem_39_1_R0_data;
  wire [7:0] R0_data_39_2 = mem_39_2_R0_data;
  wire [7:0] R0_data_39_3 = mem_39_3_R0_data;
  wire [7:0] R0_data_39_4 = mem_39_4_R0_data;
  wire [7:0] R0_data_39_5 = mem_39_5_R0_data;
  wire [7:0] R0_data_39_6 = mem_39_6_R0_data;
  wire [7:0] R0_data_39_7 = mem_39_7_R0_data;
  wire [63:0] R0_data_39 = {R0_data_39_7,R0_data_39_6,R0_data_39_5,R0_data_39_4,R0_data_39_3,R0_data_39_2,R0_data_39_1,
    R0_data_39_0};
  wire [7:0] R0_data_40_0 = mem_40_0_R0_data;
  wire [7:0] R0_data_40_1 = mem_40_1_R0_data;
  wire [7:0] R0_data_40_2 = mem_40_2_R0_data;
  wire [7:0] R0_data_40_3 = mem_40_3_R0_data;
  wire [7:0] R0_data_40_4 = mem_40_4_R0_data;
  wire [7:0] R0_data_40_5 = mem_40_5_R0_data;
  wire [7:0] R0_data_40_6 = mem_40_6_R0_data;
  wire [7:0] R0_data_40_7 = mem_40_7_R0_data;
  wire [63:0] R0_data_40 = {R0_data_40_7,R0_data_40_6,R0_data_40_5,R0_data_40_4,R0_data_40_3,R0_data_40_2,R0_data_40_1,
    R0_data_40_0};
  wire [7:0] R0_data_41_0 = mem_41_0_R0_data;
  wire [7:0] R0_data_41_1 = mem_41_1_R0_data;
  wire [7:0] R0_data_41_2 = mem_41_2_R0_data;
  wire [7:0] R0_data_41_3 = mem_41_3_R0_data;
  wire [7:0] R0_data_41_4 = mem_41_4_R0_data;
  wire [7:0] R0_data_41_5 = mem_41_5_R0_data;
  wire [7:0] R0_data_41_6 = mem_41_6_R0_data;
  wire [7:0] R0_data_41_7 = mem_41_7_R0_data;
  wire [63:0] R0_data_41 = {R0_data_41_7,R0_data_41_6,R0_data_41_5,R0_data_41_4,R0_data_41_3,R0_data_41_2,R0_data_41_1,
    R0_data_41_0};
  wire [7:0] R0_data_42_0 = mem_42_0_R0_data;
  wire [7:0] R0_data_42_1 = mem_42_1_R0_data;
  wire [7:0] R0_data_42_2 = mem_42_2_R0_data;
  wire [7:0] R0_data_42_3 = mem_42_3_R0_data;
  wire [7:0] R0_data_42_4 = mem_42_4_R0_data;
  wire [7:0] R0_data_42_5 = mem_42_5_R0_data;
  wire [7:0] R0_data_42_6 = mem_42_6_R0_data;
  wire [7:0] R0_data_42_7 = mem_42_7_R0_data;
  wire [63:0] R0_data_42 = {R0_data_42_7,R0_data_42_6,R0_data_42_5,R0_data_42_4,R0_data_42_3,R0_data_42_2,R0_data_42_1,
    R0_data_42_0};
  wire [7:0] R0_data_43_0 = mem_43_0_R0_data;
  wire [7:0] R0_data_43_1 = mem_43_1_R0_data;
  wire [7:0] R0_data_43_2 = mem_43_2_R0_data;
  wire [7:0] R0_data_43_3 = mem_43_3_R0_data;
  wire [7:0] R0_data_43_4 = mem_43_4_R0_data;
  wire [7:0] R0_data_43_5 = mem_43_5_R0_data;
  wire [7:0] R0_data_43_6 = mem_43_6_R0_data;
  wire [7:0] R0_data_43_7 = mem_43_7_R0_data;
  wire [63:0] R0_data_43 = {R0_data_43_7,R0_data_43_6,R0_data_43_5,R0_data_43_4,R0_data_43_3,R0_data_43_2,R0_data_43_1,
    R0_data_43_0};
  wire [7:0] R0_data_44_0 = mem_44_0_R0_data;
  wire [7:0] R0_data_44_1 = mem_44_1_R0_data;
  wire [7:0] R0_data_44_2 = mem_44_2_R0_data;
  wire [7:0] R0_data_44_3 = mem_44_3_R0_data;
  wire [7:0] R0_data_44_4 = mem_44_4_R0_data;
  wire [7:0] R0_data_44_5 = mem_44_5_R0_data;
  wire [7:0] R0_data_44_6 = mem_44_6_R0_data;
  wire [7:0] R0_data_44_7 = mem_44_7_R0_data;
  wire [63:0] R0_data_44 = {R0_data_44_7,R0_data_44_6,R0_data_44_5,R0_data_44_4,R0_data_44_3,R0_data_44_2,R0_data_44_1,
    R0_data_44_0};
  wire [7:0] R0_data_45_0 = mem_45_0_R0_data;
  wire [7:0] R0_data_45_1 = mem_45_1_R0_data;
  wire [7:0] R0_data_45_2 = mem_45_2_R0_data;
  wire [7:0] R0_data_45_3 = mem_45_3_R0_data;
  wire [7:0] R0_data_45_4 = mem_45_4_R0_data;
  wire [7:0] R0_data_45_5 = mem_45_5_R0_data;
  wire [7:0] R0_data_45_6 = mem_45_6_R0_data;
  wire [7:0] R0_data_45_7 = mem_45_7_R0_data;
  wire [63:0] R0_data_45 = {R0_data_45_7,R0_data_45_6,R0_data_45_5,R0_data_45_4,R0_data_45_3,R0_data_45_2,R0_data_45_1,
    R0_data_45_0};
  wire [7:0] R0_data_46_0 = mem_46_0_R0_data;
  wire [7:0] R0_data_46_1 = mem_46_1_R0_data;
  wire [7:0] R0_data_46_2 = mem_46_2_R0_data;
  wire [7:0] R0_data_46_3 = mem_46_3_R0_data;
  wire [7:0] R0_data_46_4 = mem_46_4_R0_data;
  wire [7:0] R0_data_46_5 = mem_46_5_R0_data;
  wire [7:0] R0_data_46_6 = mem_46_6_R0_data;
  wire [7:0] R0_data_46_7 = mem_46_7_R0_data;
  wire [63:0] R0_data_46 = {R0_data_46_7,R0_data_46_6,R0_data_46_5,R0_data_46_4,R0_data_46_3,R0_data_46_2,R0_data_46_1,
    R0_data_46_0};
  wire [7:0] R0_data_47_0 = mem_47_0_R0_data;
  wire [7:0] R0_data_47_1 = mem_47_1_R0_data;
  wire [7:0] R0_data_47_2 = mem_47_2_R0_data;
  wire [7:0] R0_data_47_3 = mem_47_3_R0_data;
  wire [7:0] R0_data_47_4 = mem_47_4_R0_data;
  wire [7:0] R0_data_47_5 = mem_47_5_R0_data;
  wire [7:0] R0_data_47_6 = mem_47_6_R0_data;
  wire [7:0] R0_data_47_7 = mem_47_7_R0_data;
  wire [63:0] R0_data_47 = {R0_data_47_7,R0_data_47_6,R0_data_47_5,R0_data_47_4,R0_data_47_3,R0_data_47_2,R0_data_47_1,
    R0_data_47_0};
  wire [7:0] R0_data_48_0 = mem_48_0_R0_data;
  wire [7:0] R0_data_48_1 = mem_48_1_R0_data;
  wire [7:0] R0_data_48_2 = mem_48_2_R0_data;
  wire [7:0] R0_data_48_3 = mem_48_3_R0_data;
  wire [7:0] R0_data_48_4 = mem_48_4_R0_data;
  wire [7:0] R0_data_48_5 = mem_48_5_R0_data;
  wire [7:0] R0_data_48_6 = mem_48_6_R0_data;
  wire [7:0] R0_data_48_7 = mem_48_7_R0_data;
  wire [63:0] R0_data_48 = {R0_data_48_7,R0_data_48_6,R0_data_48_5,R0_data_48_4,R0_data_48_3,R0_data_48_2,R0_data_48_1,
    R0_data_48_0};
  wire [7:0] R0_data_49_0 = mem_49_0_R0_data;
  wire [7:0] R0_data_49_1 = mem_49_1_R0_data;
  wire [7:0] R0_data_49_2 = mem_49_2_R0_data;
  wire [7:0] R0_data_49_3 = mem_49_3_R0_data;
  wire [7:0] R0_data_49_4 = mem_49_4_R0_data;
  wire [7:0] R0_data_49_5 = mem_49_5_R0_data;
  wire [7:0] R0_data_49_6 = mem_49_6_R0_data;
  wire [7:0] R0_data_49_7 = mem_49_7_R0_data;
  wire [63:0] R0_data_49 = {R0_data_49_7,R0_data_49_6,R0_data_49_5,R0_data_49_4,R0_data_49_3,R0_data_49_2,R0_data_49_1,
    R0_data_49_0};
  wire [7:0] R0_data_50_0 = mem_50_0_R0_data;
  wire [7:0] R0_data_50_1 = mem_50_1_R0_data;
  wire [7:0] R0_data_50_2 = mem_50_2_R0_data;
  wire [7:0] R0_data_50_3 = mem_50_3_R0_data;
  wire [7:0] R0_data_50_4 = mem_50_4_R0_data;
  wire [7:0] R0_data_50_5 = mem_50_5_R0_data;
  wire [7:0] R0_data_50_6 = mem_50_6_R0_data;
  wire [7:0] R0_data_50_7 = mem_50_7_R0_data;
  wire [63:0] R0_data_50 = {R0_data_50_7,R0_data_50_6,R0_data_50_5,R0_data_50_4,R0_data_50_3,R0_data_50_2,R0_data_50_1,
    R0_data_50_0};
  wire [7:0] R0_data_51_0 = mem_51_0_R0_data;
  wire [7:0] R0_data_51_1 = mem_51_1_R0_data;
  wire [7:0] R0_data_51_2 = mem_51_2_R0_data;
  wire [7:0] R0_data_51_3 = mem_51_3_R0_data;
  wire [7:0] R0_data_51_4 = mem_51_4_R0_data;
  wire [7:0] R0_data_51_5 = mem_51_5_R0_data;
  wire [7:0] R0_data_51_6 = mem_51_6_R0_data;
  wire [7:0] R0_data_51_7 = mem_51_7_R0_data;
  wire [63:0] R0_data_51 = {R0_data_51_7,R0_data_51_6,R0_data_51_5,R0_data_51_4,R0_data_51_3,R0_data_51_2,R0_data_51_1,
    R0_data_51_0};
  wire [7:0] R0_data_52_0 = mem_52_0_R0_data;
  wire [7:0] R0_data_52_1 = mem_52_1_R0_data;
  wire [7:0] R0_data_52_2 = mem_52_2_R0_data;
  wire [7:0] R0_data_52_3 = mem_52_3_R0_data;
  wire [7:0] R0_data_52_4 = mem_52_4_R0_data;
  wire [7:0] R0_data_52_5 = mem_52_5_R0_data;
  wire [7:0] R0_data_52_6 = mem_52_6_R0_data;
  wire [7:0] R0_data_52_7 = mem_52_7_R0_data;
  wire [63:0] R0_data_52 = {R0_data_52_7,R0_data_52_6,R0_data_52_5,R0_data_52_4,R0_data_52_3,R0_data_52_2,R0_data_52_1,
    R0_data_52_0};
  wire [7:0] R0_data_53_0 = mem_53_0_R0_data;
  wire [7:0] R0_data_53_1 = mem_53_1_R0_data;
  wire [7:0] R0_data_53_2 = mem_53_2_R0_data;
  wire [7:0] R0_data_53_3 = mem_53_3_R0_data;
  wire [7:0] R0_data_53_4 = mem_53_4_R0_data;
  wire [7:0] R0_data_53_5 = mem_53_5_R0_data;
  wire [7:0] R0_data_53_6 = mem_53_6_R0_data;
  wire [7:0] R0_data_53_7 = mem_53_7_R0_data;
  wire [63:0] R0_data_53 = {R0_data_53_7,R0_data_53_6,R0_data_53_5,R0_data_53_4,R0_data_53_3,R0_data_53_2,R0_data_53_1,
    R0_data_53_0};
  wire [7:0] R0_data_54_0 = mem_54_0_R0_data;
  wire [7:0] R0_data_54_1 = mem_54_1_R0_data;
  wire [7:0] R0_data_54_2 = mem_54_2_R0_data;
  wire [7:0] R0_data_54_3 = mem_54_3_R0_data;
  wire [7:0] R0_data_54_4 = mem_54_4_R0_data;
  wire [7:0] R0_data_54_5 = mem_54_5_R0_data;
  wire [7:0] R0_data_54_6 = mem_54_6_R0_data;
  wire [7:0] R0_data_54_7 = mem_54_7_R0_data;
  wire [63:0] R0_data_54 = {R0_data_54_7,R0_data_54_6,R0_data_54_5,R0_data_54_4,R0_data_54_3,R0_data_54_2,R0_data_54_1,
    R0_data_54_0};
  wire [7:0] R0_data_55_0 = mem_55_0_R0_data;
  wire [7:0] R0_data_55_1 = mem_55_1_R0_data;
  wire [7:0] R0_data_55_2 = mem_55_2_R0_data;
  wire [7:0] R0_data_55_3 = mem_55_3_R0_data;
  wire [7:0] R0_data_55_4 = mem_55_4_R0_data;
  wire [7:0] R0_data_55_5 = mem_55_5_R0_data;
  wire [7:0] R0_data_55_6 = mem_55_6_R0_data;
  wire [7:0] R0_data_55_7 = mem_55_7_R0_data;
  wire [63:0] R0_data_55 = {R0_data_55_7,R0_data_55_6,R0_data_55_5,R0_data_55_4,R0_data_55_3,R0_data_55_2,R0_data_55_1,
    R0_data_55_0};
  wire [7:0] R0_data_56_0 = mem_56_0_R0_data;
  wire [7:0] R0_data_56_1 = mem_56_1_R0_data;
  wire [7:0] R0_data_56_2 = mem_56_2_R0_data;
  wire [7:0] R0_data_56_3 = mem_56_3_R0_data;
  wire [7:0] R0_data_56_4 = mem_56_4_R0_data;
  wire [7:0] R0_data_56_5 = mem_56_5_R0_data;
  wire [7:0] R0_data_56_6 = mem_56_6_R0_data;
  wire [7:0] R0_data_56_7 = mem_56_7_R0_data;
  wire [63:0] R0_data_56 = {R0_data_56_7,R0_data_56_6,R0_data_56_5,R0_data_56_4,R0_data_56_3,R0_data_56_2,R0_data_56_1,
    R0_data_56_0};
  wire [7:0] R0_data_57_0 = mem_57_0_R0_data;
  wire [7:0] R0_data_57_1 = mem_57_1_R0_data;
  wire [7:0] R0_data_57_2 = mem_57_2_R0_data;
  wire [7:0] R0_data_57_3 = mem_57_3_R0_data;
  wire [7:0] R0_data_57_4 = mem_57_4_R0_data;
  wire [7:0] R0_data_57_5 = mem_57_5_R0_data;
  wire [7:0] R0_data_57_6 = mem_57_6_R0_data;
  wire [7:0] R0_data_57_7 = mem_57_7_R0_data;
  wire [63:0] R0_data_57 = {R0_data_57_7,R0_data_57_6,R0_data_57_5,R0_data_57_4,R0_data_57_3,R0_data_57_2,R0_data_57_1,
    R0_data_57_0};
  wire [7:0] R0_data_58_0 = mem_58_0_R0_data;
  wire [7:0] R0_data_58_1 = mem_58_1_R0_data;
  wire [7:0] R0_data_58_2 = mem_58_2_R0_data;
  wire [7:0] R0_data_58_3 = mem_58_3_R0_data;
  wire [7:0] R0_data_58_4 = mem_58_4_R0_data;
  wire [7:0] R0_data_58_5 = mem_58_5_R0_data;
  wire [7:0] R0_data_58_6 = mem_58_6_R0_data;
  wire [7:0] R0_data_58_7 = mem_58_7_R0_data;
  wire [63:0] R0_data_58 = {R0_data_58_7,R0_data_58_6,R0_data_58_5,R0_data_58_4,R0_data_58_3,R0_data_58_2,R0_data_58_1,
    R0_data_58_0};
  wire [7:0] R0_data_59_0 = mem_59_0_R0_data;
  wire [7:0] R0_data_59_1 = mem_59_1_R0_data;
  wire [7:0] R0_data_59_2 = mem_59_2_R0_data;
  wire [7:0] R0_data_59_3 = mem_59_3_R0_data;
  wire [7:0] R0_data_59_4 = mem_59_4_R0_data;
  wire [7:0] R0_data_59_5 = mem_59_5_R0_data;
  wire [7:0] R0_data_59_6 = mem_59_6_R0_data;
  wire [7:0] R0_data_59_7 = mem_59_7_R0_data;
  wire [63:0] R0_data_59 = {R0_data_59_7,R0_data_59_6,R0_data_59_5,R0_data_59_4,R0_data_59_3,R0_data_59_2,R0_data_59_1,
    R0_data_59_0};
  wire [7:0] R0_data_60_0 = mem_60_0_R0_data;
  wire [7:0] R0_data_60_1 = mem_60_1_R0_data;
  wire [7:0] R0_data_60_2 = mem_60_2_R0_data;
  wire [7:0] R0_data_60_3 = mem_60_3_R0_data;
  wire [7:0] R0_data_60_4 = mem_60_4_R0_data;
  wire [7:0] R0_data_60_5 = mem_60_5_R0_data;
  wire [7:0] R0_data_60_6 = mem_60_6_R0_data;
  wire [7:0] R0_data_60_7 = mem_60_7_R0_data;
  wire [63:0] R0_data_60 = {R0_data_60_7,R0_data_60_6,R0_data_60_5,R0_data_60_4,R0_data_60_3,R0_data_60_2,R0_data_60_1,
    R0_data_60_0};
  wire [7:0] R0_data_61_0 = mem_61_0_R0_data;
  wire [7:0] R0_data_61_1 = mem_61_1_R0_data;
  wire [7:0] R0_data_61_2 = mem_61_2_R0_data;
  wire [7:0] R0_data_61_3 = mem_61_3_R0_data;
  wire [7:0] R0_data_61_4 = mem_61_4_R0_data;
  wire [7:0] R0_data_61_5 = mem_61_5_R0_data;
  wire [7:0] R0_data_61_6 = mem_61_6_R0_data;
  wire [7:0] R0_data_61_7 = mem_61_7_R0_data;
  wire [63:0] R0_data_61 = {R0_data_61_7,R0_data_61_6,R0_data_61_5,R0_data_61_4,R0_data_61_3,R0_data_61_2,R0_data_61_1,
    R0_data_61_0};
  wire [7:0] R0_data_62_0 = mem_62_0_R0_data;
  wire [7:0] R0_data_62_1 = mem_62_1_R0_data;
  wire [7:0] R0_data_62_2 = mem_62_2_R0_data;
  wire [7:0] R0_data_62_3 = mem_62_3_R0_data;
  wire [7:0] R0_data_62_4 = mem_62_4_R0_data;
  wire [7:0] R0_data_62_5 = mem_62_5_R0_data;
  wire [7:0] R0_data_62_6 = mem_62_6_R0_data;
  wire [7:0] R0_data_62_7 = mem_62_7_R0_data;
  wire [63:0] R0_data_62 = {R0_data_62_7,R0_data_62_6,R0_data_62_5,R0_data_62_4,R0_data_62_3,R0_data_62_2,R0_data_62_1,
    R0_data_62_0};
  wire [7:0] R0_data_63_0 = mem_63_0_R0_data;
  wire [7:0] R0_data_63_1 = mem_63_1_R0_data;
  wire [7:0] R0_data_63_2 = mem_63_2_R0_data;
  wire [7:0] R0_data_63_3 = mem_63_3_R0_data;
  wire [7:0] R0_data_63_4 = mem_63_4_R0_data;
  wire [7:0] R0_data_63_5 = mem_63_5_R0_data;
  wire [7:0] R0_data_63_6 = mem_63_6_R0_data;
  wire [7:0] R0_data_63_7 = mem_63_7_R0_data;
  wire [63:0] R0_data_63 = {R0_data_63_7,R0_data_63_6,R0_data_63_5,R0_data_63_4,R0_data_63_3,R0_data_63_2,R0_data_63_1,
    R0_data_63_0};
  wire [7:0] R0_data_64_0 = mem_64_0_R0_data;
  wire [7:0] R0_data_64_1 = mem_64_1_R0_data;
  wire [7:0] R0_data_64_2 = mem_64_2_R0_data;
  wire [7:0] R0_data_64_3 = mem_64_3_R0_data;
  wire [7:0] R0_data_64_4 = mem_64_4_R0_data;
  wire [7:0] R0_data_64_5 = mem_64_5_R0_data;
  wire [7:0] R0_data_64_6 = mem_64_6_R0_data;
  wire [7:0] R0_data_64_7 = mem_64_7_R0_data;
  wire [63:0] R0_data_64 = {R0_data_64_7,R0_data_64_6,R0_data_64_5,R0_data_64_4,R0_data_64_3,R0_data_64_2,R0_data_64_1,
    R0_data_64_0};
  wire [7:0] R0_data_65_0 = mem_65_0_R0_data;
  wire [7:0] R0_data_65_1 = mem_65_1_R0_data;
  wire [7:0] R0_data_65_2 = mem_65_2_R0_data;
  wire [7:0] R0_data_65_3 = mem_65_3_R0_data;
  wire [7:0] R0_data_65_4 = mem_65_4_R0_data;
  wire [7:0] R0_data_65_5 = mem_65_5_R0_data;
  wire [7:0] R0_data_65_6 = mem_65_6_R0_data;
  wire [7:0] R0_data_65_7 = mem_65_7_R0_data;
  wire [63:0] R0_data_65 = {R0_data_65_7,R0_data_65_6,R0_data_65_5,R0_data_65_4,R0_data_65_3,R0_data_65_2,R0_data_65_1,
    R0_data_65_0};
  wire [7:0] R0_data_66_0 = mem_66_0_R0_data;
  wire [7:0] R0_data_66_1 = mem_66_1_R0_data;
  wire [7:0] R0_data_66_2 = mem_66_2_R0_data;
  wire [7:0] R0_data_66_3 = mem_66_3_R0_data;
  wire [7:0] R0_data_66_4 = mem_66_4_R0_data;
  wire [7:0] R0_data_66_5 = mem_66_5_R0_data;
  wire [7:0] R0_data_66_6 = mem_66_6_R0_data;
  wire [7:0] R0_data_66_7 = mem_66_7_R0_data;
  wire [63:0] R0_data_66 = {R0_data_66_7,R0_data_66_6,R0_data_66_5,R0_data_66_4,R0_data_66_3,R0_data_66_2,R0_data_66_1,
    R0_data_66_0};
  wire [7:0] R0_data_67_0 = mem_67_0_R0_data;
  wire [7:0] R0_data_67_1 = mem_67_1_R0_data;
  wire [7:0] R0_data_67_2 = mem_67_2_R0_data;
  wire [7:0] R0_data_67_3 = mem_67_3_R0_data;
  wire [7:0] R0_data_67_4 = mem_67_4_R0_data;
  wire [7:0] R0_data_67_5 = mem_67_5_R0_data;
  wire [7:0] R0_data_67_6 = mem_67_6_R0_data;
  wire [7:0] R0_data_67_7 = mem_67_7_R0_data;
  wire [63:0] R0_data_67 = {R0_data_67_7,R0_data_67_6,R0_data_67_5,R0_data_67_4,R0_data_67_3,R0_data_67_2,R0_data_67_1,
    R0_data_67_0};
  wire [7:0] R0_data_68_0 = mem_68_0_R0_data;
  wire [7:0] R0_data_68_1 = mem_68_1_R0_data;
  wire [7:0] R0_data_68_2 = mem_68_2_R0_data;
  wire [7:0] R0_data_68_3 = mem_68_3_R0_data;
  wire [7:0] R0_data_68_4 = mem_68_4_R0_data;
  wire [7:0] R0_data_68_5 = mem_68_5_R0_data;
  wire [7:0] R0_data_68_6 = mem_68_6_R0_data;
  wire [7:0] R0_data_68_7 = mem_68_7_R0_data;
  wire [63:0] R0_data_68 = {R0_data_68_7,R0_data_68_6,R0_data_68_5,R0_data_68_4,R0_data_68_3,R0_data_68_2,R0_data_68_1,
    R0_data_68_0};
  wire [7:0] R0_data_69_0 = mem_69_0_R0_data;
  wire [7:0] R0_data_69_1 = mem_69_1_R0_data;
  wire [7:0] R0_data_69_2 = mem_69_2_R0_data;
  wire [7:0] R0_data_69_3 = mem_69_3_R0_data;
  wire [7:0] R0_data_69_4 = mem_69_4_R0_data;
  wire [7:0] R0_data_69_5 = mem_69_5_R0_data;
  wire [7:0] R0_data_69_6 = mem_69_6_R0_data;
  wire [7:0] R0_data_69_7 = mem_69_7_R0_data;
  wire [63:0] R0_data_69 = {R0_data_69_7,R0_data_69_6,R0_data_69_5,R0_data_69_4,R0_data_69_3,R0_data_69_2,R0_data_69_1,
    R0_data_69_0};
  wire [7:0] R0_data_70_0 = mem_70_0_R0_data;
  wire [7:0] R0_data_70_1 = mem_70_1_R0_data;
  wire [7:0] R0_data_70_2 = mem_70_2_R0_data;
  wire [7:0] R0_data_70_3 = mem_70_3_R0_data;
  wire [7:0] R0_data_70_4 = mem_70_4_R0_data;
  wire [7:0] R0_data_70_5 = mem_70_5_R0_data;
  wire [7:0] R0_data_70_6 = mem_70_6_R0_data;
  wire [7:0] R0_data_70_7 = mem_70_7_R0_data;
  wire [63:0] R0_data_70 = {R0_data_70_7,R0_data_70_6,R0_data_70_5,R0_data_70_4,R0_data_70_3,R0_data_70_2,R0_data_70_1,
    R0_data_70_0};
  wire [7:0] R0_data_71_0 = mem_71_0_R0_data;
  wire [7:0] R0_data_71_1 = mem_71_1_R0_data;
  wire [7:0] R0_data_71_2 = mem_71_2_R0_data;
  wire [7:0] R0_data_71_3 = mem_71_3_R0_data;
  wire [7:0] R0_data_71_4 = mem_71_4_R0_data;
  wire [7:0] R0_data_71_5 = mem_71_5_R0_data;
  wire [7:0] R0_data_71_6 = mem_71_6_R0_data;
  wire [7:0] R0_data_71_7 = mem_71_7_R0_data;
  wire [63:0] R0_data_71 = {R0_data_71_7,R0_data_71_6,R0_data_71_5,R0_data_71_4,R0_data_71_3,R0_data_71_2,R0_data_71_1,
    R0_data_71_0};
  wire [7:0] R0_data_72_0 = mem_72_0_R0_data;
  wire [7:0] R0_data_72_1 = mem_72_1_R0_data;
  wire [7:0] R0_data_72_2 = mem_72_2_R0_data;
  wire [7:0] R0_data_72_3 = mem_72_3_R0_data;
  wire [7:0] R0_data_72_4 = mem_72_4_R0_data;
  wire [7:0] R0_data_72_5 = mem_72_5_R0_data;
  wire [7:0] R0_data_72_6 = mem_72_6_R0_data;
  wire [7:0] R0_data_72_7 = mem_72_7_R0_data;
  wire [63:0] R0_data_72 = {R0_data_72_7,R0_data_72_6,R0_data_72_5,R0_data_72_4,R0_data_72_3,R0_data_72_2,R0_data_72_1,
    R0_data_72_0};
  wire [7:0] R0_data_73_0 = mem_73_0_R0_data;
  wire [7:0] R0_data_73_1 = mem_73_1_R0_data;
  wire [7:0] R0_data_73_2 = mem_73_2_R0_data;
  wire [7:0] R0_data_73_3 = mem_73_3_R0_data;
  wire [7:0] R0_data_73_4 = mem_73_4_R0_data;
  wire [7:0] R0_data_73_5 = mem_73_5_R0_data;
  wire [7:0] R0_data_73_6 = mem_73_6_R0_data;
  wire [7:0] R0_data_73_7 = mem_73_7_R0_data;
  wire [63:0] R0_data_73 = {R0_data_73_7,R0_data_73_6,R0_data_73_5,R0_data_73_4,R0_data_73_3,R0_data_73_2,R0_data_73_1,
    R0_data_73_0};
  wire [7:0] R0_data_74_0 = mem_74_0_R0_data;
  wire [7:0] R0_data_74_1 = mem_74_1_R0_data;
  wire [7:0] R0_data_74_2 = mem_74_2_R0_data;
  wire [7:0] R0_data_74_3 = mem_74_3_R0_data;
  wire [7:0] R0_data_74_4 = mem_74_4_R0_data;
  wire [7:0] R0_data_74_5 = mem_74_5_R0_data;
  wire [7:0] R0_data_74_6 = mem_74_6_R0_data;
  wire [7:0] R0_data_74_7 = mem_74_7_R0_data;
  wire [63:0] R0_data_74 = {R0_data_74_7,R0_data_74_6,R0_data_74_5,R0_data_74_4,R0_data_74_3,R0_data_74_2,R0_data_74_1,
    R0_data_74_0};
  wire [7:0] R0_data_75_0 = mem_75_0_R0_data;
  wire [7:0] R0_data_75_1 = mem_75_1_R0_data;
  wire [7:0] R0_data_75_2 = mem_75_2_R0_data;
  wire [7:0] R0_data_75_3 = mem_75_3_R0_data;
  wire [7:0] R0_data_75_4 = mem_75_4_R0_data;
  wire [7:0] R0_data_75_5 = mem_75_5_R0_data;
  wire [7:0] R0_data_75_6 = mem_75_6_R0_data;
  wire [7:0] R0_data_75_7 = mem_75_7_R0_data;
  wire [63:0] R0_data_75 = {R0_data_75_7,R0_data_75_6,R0_data_75_5,R0_data_75_4,R0_data_75_3,R0_data_75_2,R0_data_75_1,
    R0_data_75_0};
  wire [7:0] R0_data_76_0 = mem_76_0_R0_data;
  wire [7:0] R0_data_76_1 = mem_76_1_R0_data;
  wire [7:0] R0_data_76_2 = mem_76_2_R0_data;
  wire [7:0] R0_data_76_3 = mem_76_3_R0_data;
  wire [7:0] R0_data_76_4 = mem_76_4_R0_data;
  wire [7:0] R0_data_76_5 = mem_76_5_R0_data;
  wire [7:0] R0_data_76_6 = mem_76_6_R0_data;
  wire [7:0] R0_data_76_7 = mem_76_7_R0_data;
  wire [63:0] R0_data_76 = {R0_data_76_7,R0_data_76_6,R0_data_76_5,R0_data_76_4,R0_data_76_3,R0_data_76_2,R0_data_76_1,
    R0_data_76_0};
  wire [7:0] R0_data_77_0 = mem_77_0_R0_data;
  wire [7:0] R0_data_77_1 = mem_77_1_R0_data;
  wire [7:0] R0_data_77_2 = mem_77_2_R0_data;
  wire [7:0] R0_data_77_3 = mem_77_3_R0_data;
  wire [7:0] R0_data_77_4 = mem_77_4_R0_data;
  wire [7:0] R0_data_77_5 = mem_77_5_R0_data;
  wire [7:0] R0_data_77_6 = mem_77_6_R0_data;
  wire [7:0] R0_data_77_7 = mem_77_7_R0_data;
  wire [63:0] R0_data_77 = {R0_data_77_7,R0_data_77_6,R0_data_77_5,R0_data_77_4,R0_data_77_3,R0_data_77_2,R0_data_77_1,
    R0_data_77_0};
  wire [7:0] R0_data_78_0 = mem_78_0_R0_data;
  wire [7:0] R0_data_78_1 = mem_78_1_R0_data;
  wire [7:0] R0_data_78_2 = mem_78_2_R0_data;
  wire [7:0] R0_data_78_3 = mem_78_3_R0_data;
  wire [7:0] R0_data_78_4 = mem_78_4_R0_data;
  wire [7:0] R0_data_78_5 = mem_78_5_R0_data;
  wire [7:0] R0_data_78_6 = mem_78_6_R0_data;
  wire [7:0] R0_data_78_7 = mem_78_7_R0_data;
  wire [63:0] R0_data_78 = {R0_data_78_7,R0_data_78_6,R0_data_78_5,R0_data_78_4,R0_data_78_3,R0_data_78_2,R0_data_78_1,
    R0_data_78_0};
  wire [7:0] R0_data_79_0 = mem_79_0_R0_data;
  wire [7:0] R0_data_79_1 = mem_79_1_R0_data;
  wire [7:0] R0_data_79_2 = mem_79_2_R0_data;
  wire [7:0] R0_data_79_3 = mem_79_3_R0_data;
  wire [7:0] R0_data_79_4 = mem_79_4_R0_data;
  wire [7:0] R0_data_79_5 = mem_79_5_R0_data;
  wire [7:0] R0_data_79_6 = mem_79_6_R0_data;
  wire [7:0] R0_data_79_7 = mem_79_7_R0_data;
  wire [63:0] R0_data_79 = {R0_data_79_7,R0_data_79_6,R0_data_79_5,R0_data_79_4,R0_data_79_3,R0_data_79_2,R0_data_79_1,
    R0_data_79_0};
  wire [7:0] R0_data_80_0 = mem_80_0_R0_data;
  wire [7:0] R0_data_80_1 = mem_80_1_R0_data;
  wire [7:0] R0_data_80_2 = mem_80_2_R0_data;
  wire [7:0] R0_data_80_3 = mem_80_3_R0_data;
  wire [7:0] R0_data_80_4 = mem_80_4_R0_data;
  wire [7:0] R0_data_80_5 = mem_80_5_R0_data;
  wire [7:0] R0_data_80_6 = mem_80_6_R0_data;
  wire [7:0] R0_data_80_7 = mem_80_7_R0_data;
  wire [63:0] R0_data_80 = {R0_data_80_7,R0_data_80_6,R0_data_80_5,R0_data_80_4,R0_data_80_3,R0_data_80_2,R0_data_80_1,
    R0_data_80_0};
  wire [7:0] R0_data_81_0 = mem_81_0_R0_data;
  wire [7:0] R0_data_81_1 = mem_81_1_R0_data;
  wire [7:0] R0_data_81_2 = mem_81_2_R0_data;
  wire [7:0] R0_data_81_3 = mem_81_3_R0_data;
  wire [7:0] R0_data_81_4 = mem_81_4_R0_data;
  wire [7:0] R0_data_81_5 = mem_81_5_R0_data;
  wire [7:0] R0_data_81_6 = mem_81_6_R0_data;
  wire [7:0] R0_data_81_7 = mem_81_7_R0_data;
  wire [63:0] R0_data_81 = {R0_data_81_7,R0_data_81_6,R0_data_81_5,R0_data_81_4,R0_data_81_3,R0_data_81_2,R0_data_81_1,
    R0_data_81_0};
  wire [7:0] R0_data_82_0 = mem_82_0_R0_data;
  wire [7:0] R0_data_82_1 = mem_82_1_R0_data;
  wire [7:0] R0_data_82_2 = mem_82_2_R0_data;
  wire [7:0] R0_data_82_3 = mem_82_3_R0_data;
  wire [7:0] R0_data_82_4 = mem_82_4_R0_data;
  wire [7:0] R0_data_82_5 = mem_82_5_R0_data;
  wire [7:0] R0_data_82_6 = mem_82_6_R0_data;
  wire [7:0] R0_data_82_7 = mem_82_7_R0_data;
  wire [63:0] R0_data_82 = {R0_data_82_7,R0_data_82_6,R0_data_82_5,R0_data_82_4,R0_data_82_3,R0_data_82_2,R0_data_82_1,
    R0_data_82_0};
  wire [7:0] R0_data_83_0 = mem_83_0_R0_data;
  wire [7:0] R0_data_83_1 = mem_83_1_R0_data;
  wire [7:0] R0_data_83_2 = mem_83_2_R0_data;
  wire [7:0] R0_data_83_3 = mem_83_3_R0_data;
  wire [7:0] R0_data_83_4 = mem_83_4_R0_data;
  wire [7:0] R0_data_83_5 = mem_83_5_R0_data;
  wire [7:0] R0_data_83_6 = mem_83_6_R0_data;
  wire [7:0] R0_data_83_7 = mem_83_7_R0_data;
  wire [63:0] R0_data_83 = {R0_data_83_7,R0_data_83_6,R0_data_83_5,R0_data_83_4,R0_data_83_3,R0_data_83_2,R0_data_83_1,
    R0_data_83_0};
  wire [7:0] R0_data_84_0 = mem_84_0_R0_data;
  wire [7:0] R0_data_84_1 = mem_84_1_R0_data;
  wire [7:0] R0_data_84_2 = mem_84_2_R0_data;
  wire [7:0] R0_data_84_3 = mem_84_3_R0_data;
  wire [7:0] R0_data_84_4 = mem_84_4_R0_data;
  wire [7:0] R0_data_84_5 = mem_84_5_R0_data;
  wire [7:0] R0_data_84_6 = mem_84_6_R0_data;
  wire [7:0] R0_data_84_7 = mem_84_7_R0_data;
  wire [63:0] R0_data_84 = {R0_data_84_7,R0_data_84_6,R0_data_84_5,R0_data_84_4,R0_data_84_3,R0_data_84_2,R0_data_84_1,
    R0_data_84_0};
  wire [7:0] R0_data_85_0 = mem_85_0_R0_data;
  wire [7:0] R0_data_85_1 = mem_85_1_R0_data;
  wire [7:0] R0_data_85_2 = mem_85_2_R0_data;
  wire [7:0] R0_data_85_3 = mem_85_3_R0_data;
  wire [7:0] R0_data_85_4 = mem_85_4_R0_data;
  wire [7:0] R0_data_85_5 = mem_85_5_R0_data;
  wire [7:0] R0_data_85_6 = mem_85_6_R0_data;
  wire [7:0] R0_data_85_7 = mem_85_7_R0_data;
  wire [63:0] R0_data_85 = {R0_data_85_7,R0_data_85_6,R0_data_85_5,R0_data_85_4,R0_data_85_3,R0_data_85_2,R0_data_85_1,
    R0_data_85_0};
  wire [7:0] R0_data_86_0 = mem_86_0_R0_data;
  wire [7:0] R0_data_86_1 = mem_86_1_R0_data;
  wire [7:0] R0_data_86_2 = mem_86_2_R0_data;
  wire [7:0] R0_data_86_3 = mem_86_3_R0_data;
  wire [7:0] R0_data_86_4 = mem_86_4_R0_data;
  wire [7:0] R0_data_86_5 = mem_86_5_R0_data;
  wire [7:0] R0_data_86_6 = mem_86_6_R0_data;
  wire [7:0] R0_data_86_7 = mem_86_7_R0_data;
  wire [63:0] R0_data_86 = {R0_data_86_7,R0_data_86_6,R0_data_86_5,R0_data_86_4,R0_data_86_3,R0_data_86_2,R0_data_86_1,
    R0_data_86_0};
  wire [7:0] R0_data_87_0 = mem_87_0_R0_data;
  wire [7:0] R0_data_87_1 = mem_87_1_R0_data;
  wire [7:0] R0_data_87_2 = mem_87_2_R0_data;
  wire [7:0] R0_data_87_3 = mem_87_3_R0_data;
  wire [7:0] R0_data_87_4 = mem_87_4_R0_data;
  wire [7:0] R0_data_87_5 = mem_87_5_R0_data;
  wire [7:0] R0_data_87_6 = mem_87_6_R0_data;
  wire [7:0] R0_data_87_7 = mem_87_7_R0_data;
  wire [63:0] R0_data_87 = {R0_data_87_7,R0_data_87_6,R0_data_87_5,R0_data_87_4,R0_data_87_3,R0_data_87_2,R0_data_87_1,
    R0_data_87_0};
  wire [7:0] R0_data_88_0 = mem_88_0_R0_data;
  wire [7:0] R0_data_88_1 = mem_88_1_R0_data;
  wire [7:0] R0_data_88_2 = mem_88_2_R0_data;
  wire [7:0] R0_data_88_3 = mem_88_3_R0_data;
  wire [7:0] R0_data_88_4 = mem_88_4_R0_data;
  wire [7:0] R0_data_88_5 = mem_88_5_R0_data;
  wire [7:0] R0_data_88_6 = mem_88_6_R0_data;
  wire [7:0] R0_data_88_7 = mem_88_7_R0_data;
  wire [63:0] R0_data_88 = {R0_data_88_7,R0_data_88_6,R0_data_88_5,R0_data_88_4,R0_data_88_3,R0_data_88_2,R0_data_88_1,
    R0_data_88_0};
  wire [7:0] R0_data_89_0 = mem_89_0_R0_data;
  wire [7:0] R0_data_89_1 = mem_89_1_R0_data;
  wire [7:0] R0_data_89_2 = mem_89_2_R0_data;
  wire [7:0] R0_data_89_3 = mem_89_3_R0_data;
  wire [7:0] R0_data_89_4 = mem_89_4_R0_data;
  wire [7:0] R0_data_89_5 = mem_89_5_R0_data;
  wire [7:0] R0_data_89_6 = mem_89_6_R0_data;
  wire [7:0] R0_data_89_7 = mem_89_7_R0_data;
  wire [63:0] R0_data_89 = {R0_data_89_7,R0_data_89_6,R0_data_89_5,R0_data_89_4,R0_data_89_3,R0_data_89_2,R0_data_89_1,
    R0_data_89_0};
  wire [7:0] R0_data_90_0 = mem_90_0_R0_data;
  wire [7:0] R0_data_90_1 = mem_90_1_R0_data;
  wire [7:0] R0_data_90_2 = mem_90_2_R0_data;
  wire [7:0] R0_data_90_3 = mem_90_3_R0_data;
  wire [7:0] R0_data_90_4 = mem_90_4_R0_data;
  wire [7:0] R0_data_90_5 = mem_90_5_R0_data;
  wire [7:0] R0_data_90_6 = mem_90_6_R0_data;
  wire [7:0] R0_data_90_7 = mem_90_7_R0_data;
  wire [63:0] R0_data_90 = {R0_data_90_7,R0_data_90_6,R0_data_90_5,R0_data_90_4,R0_data_90_3,R0_data_90_2,R0_data_90_1,
    R0_data_90_0};
  wire [7:0] R0_data_91_0 = mem_91_0_R0_data;
  wire [7:0] R0_data_91_1 = mem_91_1_R0_data;
  wire [7:0] R0_data_91_2 = mem_91_2_R0_data;
  wire [7:0] R0_data_91_3 = mem_91_3_R0_data;
  wire [7:0] R0_data_91_4 = mem_91_4_R0_data;
  wire [7:0] R0_data_91_5 = mem_91_5_R0_data;
  wire [7:0] R0_data_91_6 = mem_91_6_R0_data;
  wire [7:0] R0_data_91_7 = mem_91_7_R0_data;
  wire [63:0] R0_data_91 = {R0_data_91_7,R0_data_91_6,R0_data_91_5,R0_data_91_4,R0_data_91_3,R0_data_91_2,R0_data_91_1,
    R0_data_91_0};
  wire [7:0] R0_data_92_0 = mem_92_0_R0_data;
  wire [7:0] R0_data_92_1 = mem_92_1_R0_data;
  wire [7:0] R0_data_92_2 = mem_92_2_R0_data;
  wire [7:0] R0_data_92_3 = mem_92_3_R0_data;
  wire [7:0] R0_data_92_4 = mem_92_4_R0_data;
  wire [7:0] R0_data_92_5 = mem_92_5_R0_data;
  wire [7:0] R0_data_92_6 = mem_92_6_R0_data;
  wire [7:0] R0_data_92_7 = mem_92_7_R0_data;
  wire [63:0] R0_data_92 = {R0_data_92_7,R0_data_92_6,R0_data_92_5,R0_data_92_4,R0_data_92_3,R0_data_92_2,R0_data_92_1,
    R0_data_92_0};
  wire [7:0] R0_data_93_0 = mem_93_0_R0_data;
  wire [7:0] R0_data_93_1 = mem_93_1_R0_data;
  wire [7:0] R0_data_93_2 = mem_93_2_R0_data;
  wire [7:0] R0_data_93_3 = mem_93_3_R0_data;
  wire [7:0] R0_data_93_4 = mem_93_4_R0_data;
  wire [7:0] R0_data_93_5 = mem_93_5_R0_data;
  wire [7:0] R0_data_93_6 = mem_93_6_R0_data;
  wire [7:0] R0_data_93_7 = mem_93_7_R0_data;
  wire [63:0] R0_data_93 = {R0_data_93_7,R0_data_93_6,R0_data_93_5,R0_data_93_4,R0_data_93_3,R0_data_93_2,R0_data_93_1,
    R0_data_93_0};
  wire [7:0] R0_data_94_0 = mem_94_0_R0_data;
  wire [7:0] R0_data_94_1 = mem_94_1_R0_data;
  wire [7:0] R0_data_94_2 = mem_94_2_R0_data;
  wire [7:0] R0_data_94_3 = mem_94_3_R0_data;
  wire [7:0] R0_data_94_4 = mem_94_4_R0_data;
  wire [7:0] R0_data_94_5 = mem_94_5_R0_data;
  wire [7:0] R0_data_94_6 = mem_94_6_R0_data;
  wire [7:0] R0_data_94_7 = mem_94_7_R0_data;
  wire [63:0] R0_data_94 = {R0_data_94_7,R0_data_94_6,R0_data_94_5,R0_data_94_4,R0_data_94_3,R0_data_94_2,R0_data_94_1,
    R0_data_94_0};
  wire [7:0] R0_data_95_0 = mem_95_0_R0_data;
  wire [7:0] R0_data_95_1 = mem_95_1_R0_data;
  wire [7:0] R0_data_95_2 = mem_95_2_R0_data;
  wire [7:0] R0_data_95_3 = mem_95_3_R0_data;
  wire [7:0] R0_data_95_4 = mem_95_4_R0_data;
  wire [7:0] R0_data_95_5 = mem_95_5_R0_data;
  wire [7:0] R0_data_95_6 = mem_95_6_R0_data;
  wire [7:0] R0_data_95_7 = mem_95_7_R0_data;
  wire [63:0] R0_data_95 = {R0_data_95_7,R0_data_95_6,R0_data_95_5,R0_data_95_4,R0_data_95_3,R0_data_95_2,R0_data_95_1,
    R0_data_95_0};
  wire [7:0] R0_data_96_0 = mem_96_0_R0_data;
  wire [7:0] R0_data_96_1 = mem_96_1_R0_data;
  wire [7:0] R0_data_96_2 = mem_96_2_R0_data;
  wire [7:0] R0_data_96_3 = mem_96_3_R0_data;
  wire [7:0] R0_data_96_4 = mem_96_4_R0_data;
  wire [7:0] R0_data_96_5 = mem_96_5_R0_data;
  wire [7:0] R0_data_96_6 = mem_96_6_R0_data;
  wire [7:0] R0_data_96_7 = mem_96_7_R0_data;
  wire [63:0] R0_data_96 = {R0_data_96_7,R0_data_96_6,R0_data_96_5,R0_data_96_4,R0_data_96_3,R0_data_96_2,R0_data_96_1,
    R0_data_96_0};
  wire [7:0] R0_data_97_0 = mem_97_0_R0_data;
  wire [7:0] R0_data_97_1 = mem_97_1_R0_data;
  wire [7:0] R0_data_97_2 = mem_97_2_R0_data;
  wire [7:0] R0_data_97_3 = mem_97_3_R0_data;
  wire [7:0] R0_data_97_4 = mem_97_4_R0_data;
  wire [7:0] R0_data_97_5 = mem_97_5_R0_data;
  wire [7:0] R0_data_97_6 = mem_97_6_R0_data;
  wire [7:0] R0_data_97_7 = mem_97_7_R0_data;
  wire [63:0] R0_data_97 = {R0_data_97_7,R0_data_97_6,R0_data_97_5,R0_data_97_4,R0_data_97_3,R0_data_97_2,R0_data_97_1,
    R0_data_97_0};
  wire [7:0] R0_data_98_0 = mem_98_0_R0_data;
  wire [7:0] R0_data_98_1 = mem_98_1_R0_data;
  wire [7:0] R0_data_98_2 = mem_98_2_R0_data;
  wire [7:0] R0_data_98_3 = mem_98_3_R0_data;
  wire [7:0] R0_data_98_4 = mem_98_4_R0_data;
  wire [7:0] R0_data_98_5 = mem_98_5_R0_data;
  wire [7:0] R0_data_98_6 = mem_98_6_R0_data;
  wire [7:0] R0_data_98_7 = mem_98_7_R0_data;
  wire [63:0] R0_data_98 = {R0_data_98_7,R0_data_98_6,R0_data_98_5,R0_data_98_4,R0_data_98_3,R0_data_98_2,R0_data_98_1,
    R0_data_98_0};
  wire [7:0] R0_data_99_0 = mem_99_0_R0_data;
  wire [7:0] R0_data_99_1 = mem_99_1_R0_data;
  wire [7:0] R0_data_99_2 = mem_99_2_R0_data;
  wire [7:0] R0_data_99_3 = mem_99_3_R0_data;
  wire [7:0] R0_data_99_4 = mem_99_4_R0_data;
  wire [7:0] R0_data_99_5 = mem_99_5_R0_data;
  wire [7:0] R0_data_99_6 = mem_99_6_R0_data;
  wire [7:0] R0_data_99_7 = mem_99_7_R0_data;
  wire [63:0] R0_data_99 = {R0_data_99_7,R0_data_99_6,R0_data_99_5,R0_data_99_4,R0_data_99_3,R0_data_99_2,R0_data_99_1,
    R0_data_99_0};
  wire [7:0] R0_data_100_0 = mem_100_0_R0_data;
  wire [7:0] R0_data_100_1 = mem_100_1_R0_data;
  wire [7:0] R0_data_100_2 = mem_100_2_R0_data;
  wire [7:0] R0_data_100_3 = mem_100_3_R0_data;
  wire [7:0] R0_data_100_4 = mem_100_4_R0_data;
  wire [7:0] R0_data_100_5 = mem_100_5_R0_data;
  wire [7:0] R0_data_100_6 = mem_100_6_R0_data;
  wire [7:0] R0_data_100_7 = mem_100_7_R0_data;
  wire [63:0] R0_data_100 = {R0_data_100_7,R0_data_100_6,R0_data_100_5,R0_data_100_4,R0_data_100_3,R0_data_100_2,
    R0_data_100_1,R0_data_100_0};
  wire [7:0] R0_data_101_0 = mem_101_0_R0_data;
  wire [7:0] R0_data_101_1 = mem_101_1_R0_data;
  wire [7:0] R0_data_101_2 = mem_101_2_R0_data;
  wire [7:0] R0_data_101_3 = mem_101_3_R0_data;
  wire [7:0] R0_data_101_4 = mem_101_4_R0_data;
  wire [7:0] R0_data_101_5 = mem_101_5_R0_data;
  wire [7:0] R0_data_101_6 = mem_101_6_R0_data;
  wire [7:0] R0_data_101_7 = mem_101_7_R0_data;
  wire [63:0] R0_data_101 = {R0_data_101_7,R0_data_101_6,R0_data_101_5,R0_data_101_4,R0_data_101_3,R0_data_101_2,
    R0_data_101_1,R0_data_101_0};
  wire [7:0] R0_data_102_0 = mem_102_0_R0_data;
  wire [7:0] R0_data_102_1 = mem_102_1_R0_data;
  wire [7:0] R0_data_102_2 = mem_102_2_R0_data;
  wire [7:0] R0_data_102_3 = mem_102_3_R0_data;
  wire [7:0] R0_data_102_4 = mem_102_4_R0_data;
  wire [7:0] R0_data_102_5 = mem_102_5_R0_data;
  wire [7:0] R0_data_102_6 = mem_102_6_R0_data;
  wire [7:0] R0_data_102_7 = mem_102_7_R0_data;
  wire [63:0] R0_data_102 = {R0_data_102_7,R0_data_102_6,R0_data_102_5,R0_data_102_4,R0_data_102_3,R0_data_102_2,
    R0_data_102_1,R0_data_102_0};
  wire [7:0] R0_data_103_0 = mem_103_0_R0_data;
  wire [7:0] R0_data_103_1 = mem_103_1_R0_data;
  wire [7:0] R0_data_103_2 = mem_103_2_R0_data;
  wire [7:0] R0_data_103_3 = mem_103_3_R0_data;
  wire [7:0] R0_data_103_4 = mem_103_4_R0_data;
  wire [7:0] R0_data_103_5 = mem_103_5_R0_data;
  wire [7:0] R0_data_103_6 = mem_103_6_R0_data;
  wire [7:0] R0_data_103_7 = mem_103_7_R0_data;
  wire [63:0] R0_data_103 = {R0_data_103_7,R0_data_103_6,R0_data_103_5,R0_data_103_4,R0_data_103_3,R0_data_103_2,
    R0_data_103_1,R0_data_103_0};
  wire [7:0] R0_data_104_0 = mem_104_0_R0_data;
  wire [7:0] R0_data_104_1 = mem_104_1_R0_data;
  wire [7:0] R0_data_104_2 = mem_104_2_R0_data;
  wire [7:0] R0_data_104_3 = mem_104_3_R0_data;
  wire [7:0] R0_data_104_4 = mem_104_4_R0_data;
  wire [7:0] R0_data_104_5 = mem_104_5_R0_data;
  wire [7:0] R0_data_104_6 = mem_104_6_R0_data;
  wire [7:0] R0_data_104_7 = mem_104_7_R0_data;
  wire [63:0] R0_data_104 = {R0_data_104_7,R0_data_104_6,R0_data_104_5,R0_data_104_4,R0_data_104_3,R0_data_104_2,
    R0_data_104_1,R0_data_104_0};
  wire [7:0] R0_data_105_0 = mem_105_0_R0_data;
  wire [7:0] R0_data_105_1 = mem_105_1_R0_data;
  wire [7:0] R0_data_105_2 = mem_105_2_R0_data;
  wire [7:0] R0_data_105_3 = mem_105_3_R0_data;
  wire [7:0] R0_data_105_4 = mem_105_4_R0_data;
  wire [7:0] R0_data_105_5 = mem_105_5_R0_data;
  wire [7:0] R0_data_105_6 = mem_105_6_R0_data;
  wire [7:0] R0_data_105_7 = mem_105_7_R0_data;
  wire [63:0] R0_data_105 = {R0_data_105_7,R0_data_105_6,R0_data_105_5,R0_data_105_4,R0_data_105_3,R0_data_105_2,
    R0_data_105_1,R0_data_105_0};
  wire [7:0] R0_data_106_0 = mem_106_0_R0_data;
  wire [7:0] R0_data_106_1 = mem_106_1_R0_data;
  wire [7:0] R0_data_106_2 = mem_106_2_R0_data;
  wire [7:0] R0_data_106_3 = mem_106_3_R0_data;
  wire [7:0] R0_data_106_4 = mem_106_4_R0_data;
  wire [7:0] R0_data_106_5 = mem_106_5_R0_data;
  wire [7:0] R0_data_106_6 = mem_106_6_R0_data;
  wire [7:0] R0_data_106_7 = mem_106_7_R0_data;
  wire [63:0] R0_data_106 = {R0_data_106_7,R0_data_106_6,R0_data_106_5,R0_data_106_4,R0_data_106_3,R0_data_106_2,
    R0_data_106_1,R0_data_106_0};
  wire [7:0] R0_data_107_0 = mem_107_0_R0_data;
  wire [7:0] R0_data_107_1 = mem_107_1_R0_data;
  wire [7:0] R0_data_107_2 = mem_107_2_R0_data;
  wire [7:0] R0_data_107_3 = mem_107_3_R0_data;
  wire [7:0] R0_data_107_4 = mem_107_4_R0_data;
  wire [7:0] R0_data_107_5 = mem_107_5_R0_data;
  wire [7:0] R0_data_107_6 = mem_107_6_R0_data;
  wire [7:0] R0_data_107_7 = mem_107_7_R0_data;
  wire [63:0] R0_data_107 = {R0_data_107_7,R0_data_107_6,R0_data_107_5,R0_data_107_4,R0_data_107_3,R0_data_107_2,
    R0_data_107_1,R0_data_107_0};
  wire [7:0] R0_data_108_0 = mem_108_0_R0_data;
  wire [7:0] R0_data_108_1 = mem_108_1_R0_data;
  wire [7:0] R0_data_108_2 = mem_108_2_R0_data;
  wire [7:0] R0_data_108_3 = mem_108_3_R0_data;
  wire [7:0] R0_data_108_4 = mem_108_4_R0_data;
  wire [7:0] R0_data_108_5 = mem_108_5_R0_data;
  wire [7:0] R0_data_108_6 = mem_108_6_R0_data;
  wire [7:0] R0_data_108_7 = mem_108_7_R0_data;
  wire [63:0] R0_data_108 = {R0_data_108_7,R0_data_108_6,R0_data_108_5,R0_data_108_4,R0_data_108_3,R0_data_108_2,
    R0_data_108_1,R0_data_108_0};
  wire [7:0] R0_data_109_0 = mem_109_0_R0_data;
  wire [7:0] R0_data_109_1 = mem_109_1_R0_data;
  wire [7:0] R0_data_109_2 = mem_109_2_R0_data;
  wire [7:0] R0_data_109_3 = mem_109_3_R0_data;
  wire [7:0] R0_data_109_4 = mem_109_4_R0_data;
  wire [7:0] R0_data_109_5 = mem_109_5_R0_data;
  wire [7:0] R0_data_109_6 = mem_109_6_R0_data;
  wire [7:0] R0_data_109_7 = mem_109_7_R0_data;
  wire [63:0] R0_data_109 = {R0_data_109_7,R0_data_109_6,R0_data_109_5,R0_data_109_4,R0_data_109_3,R0_data_109_2,
    R0_data_109_1,R0_data_109_0};
  wire [7:0] R0_data_110_0 = mem_110_0_R0_data;
  wire [7:0] R0_data_110_1 = mem_110_1_R0_data;
  wire [7:0] R0_data_110_2 = mem_110_2_R0_data;
  wire [7:0] R0_data_110_3 = mem_110_3_R0_data;
  wire [7:0] R0_data_110_4 = mem_110_4_R0_data;
  wire [7:0] R0_data_110_5 = mem_110_5_R0_data;
  wire [7:0] R0_data_110_6 = mem_110_6_R0_data;
  wire [7:0] R0_data_110_7 = mem_110_7_R0_data;
  wire [63:0] R0_data_110 = {R0_data_110_7,R0_data_110_6,R0_data_110_5,R0_data_110_4,R0_data_110_3,R0_data_110_2,
    R0_data_110_1,R0_data_110_0};
  wire [7:0] R0_data_111_0 = mem_111_0_R0_data;
  wire [7:0] R0_data_111_1 = mem_111_1_R0_data;
  wire [7:0] R0_data_111_2 = mem_111_2_R0_data;
  wire [7:0] R0_data_111_3 = mem_111_3_R0_data;
  wire [7:0] R0_data_111_4 = mem_111_4_R0_data;
  wire [7:0] R0_data_111_5 = mem_111_5_R0_data;
  wire [7:0] R0_data_111_6 = mem_111_6_R0_data;
  wire [7:0] R0_data_111_7 = mem_111_7_R0_data;
  wire [63:0] R0_data_111 = {R0_data_111_7,R0_data_111_6,R0_data_111_5,R0_data_111_4,R0_data_111_3,R0_data_111_2,
    R0_data_111_1,R0_data_111_0};
  wire [7:0] R0_data_112_0 = mem_112_0_R0_data;
  wire [7:0] R0_data_112_1 = mem_112_1_R0_data;
  wire [7:0] R0_data_112_2 = mem_112_2_R0_data;
  wire [7:0] R0_data_112_3 = mem_112_3_R0_data;
  wire [7:0] R0_data_112_4 = mem_112_4_R0_data;
  wire [7:0] R0_data_112_5 = mem_112_5_R0_data;
  wire [7:0] R0_data_112_6 = mem_112_6_R0_data;
  wire [7:0] R0_data_112_7 = mem_112_7_R0_data;
  wire [63:0] R0_data_112 = {R0_data_112_7,R0_data_112_6,R0_data_112_5,R0_data_112_4,R0_data_112_3,R0_data_112_2,
    R0_data_112_1,R0_data_112_0};
  wire [7:0] R0_data_113_0 = mem_113_0_R0_data;
  wire [7:0] R0_data_113_1 = mem_113_1_R0_data;
  wire [7:0] R0_data_113_2 = mem_113_2_R0_data;
  wire [7:0] R0_data_113_3 = mem_113_3_R0_data;
  wire [7:0] R0_data_113_4 = mem_113_4_R0_data;
  wire [7:0] R0_data_113_5 = mem_113_5_R0_data;
  wire [7:0] R0_data_113_6 = mem_113_6_R0_data;
  wire [7:0] R0_data_113_7 = mem_113_7_R0_data;
  wire [63:0] R0_data_113 = {R0_data_113_7,R0_data_113_6,R0_data_113_5,R0_data_113_4,R0_data_113_3,R0_data_113_2,
    R0_data_113_1,R0_data_113_0};
  wire [7:0] R0_data_114_0 = mem_114_0_R0_data;
  wire [7:0] R0_data_114_1 = mem_114_1_R0_data;
  wire [7:0] R0_data_114_2 = mem_114_2_R0_data;
  wire [7:0] R0_data_114_3 = mem_114_3_R0_data;
  wire [7:0] R0_data_114_4 = mem_114_4_R0_data;
  wire [7:0] R0_data_114_5 = mem_114_5_R0_data;
  wire [7:0] R0_data_114_6 = mem_114_6_R0_data;
  wire [7:0] R0_data_114_7 = mem_114_7_R0_data;
  wire [63:0] R0_data_114 = {R0_data_114_7,R0_data_114_6,R0_data_114_5,R0_data_114_4,R0_data_114_3,R0_data_114_2,
    R0_data_114_1,R0_data_114_0};
  wire [7:0] R0_data_115_0 = mem_115_0_R0_data;
  wire [7:0] R0_data_115_1 = mem_115_1_R0_data;
  wire [7:0] R0_data_115_2 = mem_115_2_R0_data;
  wire [7:0] R0_data_115_3 = mem_115_3_R0_data;
  wire [7:0] R0_data_115_4 = mem_115_4_R0_data;
  wire [7:0] R0_data_115_5 = mem_115_5_R0_data;
  wire [7:0] R0_data_115_6 = mem_115_6_R0_data;
  wire [7:0] R0_data_115_7 = mem_115_7_R0_data;
  wire [63:0] R0_data_115 = {R0_data_115_7,R0_data_115_6,R0_data_115_5,R0_data_115_4,R0_data_115_3,R0_data_115_2,
    R0_data_115_1,R0_data_115_0};
  wire [7:0] R0_data_116_0 = mem_116_0_R0_data;
  wire [7:0] R0_data_116_1 = mem_116_1_R0_data;
  wire [7:0] R0_data_116_2 = mem_116_2_R0_data;
  wire [7:0] R0_data_116_3 = mem_116_3_R0_data;
  wire [7:0] R0_data_116_4 = mem_116_4_R0_data;
  wire [7:0] R0_data_116_5 = mem_116_5_R0_data;
  wire [7:0] R0_data_116_6 = mem_116_6_R0_data;
  wire [7:0] R0_data_116_7 = mem_116_7_R0_data;
  wire [63:0] R0_data_116 = {R0_data_116_7,R0_data_116_6,R0_data_116_5,R0_data_116_4,R0_data_116_3,R0_data_116_2,
    R0_data_116_1,R0_data_116_0};
  wire [7:0] R0_data_117_0 = mem_117_0_R0_data;
  wire [7:0] R0_data_117_1 = mem_117_1_R0_data;
  wire [7:0] R0_data_117_2 = mem_117_2_R0_data;
  wire [7:0] R0_data_117_3 = mem_117_3_R0_data;
  wire [7:0] R0_data_117_4 = mem_117_4_R0_data;
  wire [7:0] R0_data_117_5 = mem_117_5_R0_data;
  wire [7:0] R0_data_117_6 = mem_117_6_R0_data;
  wire [7:0] R0_data_117_7 = mem_117_7_R0_data;
  wire [63:0] R0_data_117 = {R0_data_117_7,R0_data_117_6,R0_data_117_5,R0_data_117_4,R0_data_117_3,R0_data_117_2,
    R0_data_117_1,R0_data_117_0};
  wire [7:0] R0_data_118_0 = mem_118_0_R0_data;
  wire [7:0] R0_data_118_1 = mem_118_1_R0_data;
  wire [7:0] R0_data_118_2 = mem_118_2_R0_data;
  wire [7:0] R0_data_118_3 = mem_118_3_R0_data;
  wire [7:0] R0_data_118_4 = mem_118_4_R0_data;
  wire [7:0] R0_data_118_5 = mem_118_5_R0_data;
  wire [7:0] R0_data_118_6 = mem_118_6_R0_data;
  wire [7:0] R0_data_118_7 = mem_118_7_R0_data;
  wire [63:0] R0_data_118 = {R0_data_118_7,R0_data_118_6,R0_data_118_5,R0_data_118_4,R0_data_118_3,R0_data_118_2,
    R0_data_118_1,R0_data_118_0};
  wire [7:0] R0_data_119_0 = mem_119_0_R0_data;
  wire [7:0] R0_data_119_1 = mem_119_1_R0_data;
  wire [7:0] R0_data_119_2 = mem_119_2_R0_data;
  wire [7:0] R0_data_119_3 = mem_119_3_R0_data;
  wire [7:0] R0_data_119_4 = mem_119_4_R0_data;
  wire [7:0] R0_data_119_5 = mem_119_5_R0_data;
  wire [7:0] R0_data_119_6 = mem_119_6_R0_data;
  wire [7:0] R0_data_119_7 = mem_119_7_R0_data;
  wire [63:0] R0_data_119 = {R0_data_119_7,R0_data_119_6,R0_data_119_5,R0_data_119_4,R0_data_119_3,R0_data_119_2,
    R0_data_119_1,R0_data_119_0};
  wire [7:0] R0_data_120_0 = mem_120_0_R0_data;
  wire [7:0] R0_data_120_1 = mem_120_1_R0_data;
  wire [7:0] R0_data_120_2 = mem_120_2_R0_data;
  wire [7:0] R0_data_120_3 = mem_120_3_R0_data;
  wire [7:0] R0_data_120_4 = mem_120_4_R0_data;
  wire [7:0] R0_data_120_5 = mem_120_5_R0_data;
  wire [7:0] R0_data_120_6 = mem_120_6_R0_data;
  wire [7:0] R0_data_120_7 = mem_120_7_R0_data;
  wire [63:0] R0_data_120 = {R0_data_120_7,R0_data_120_6,R0_data_120_5,R0_data_120_4,R0_data_120_3,R0_data_120_2,
    R0_data_120_1,R0_data_120_0};
  wire [7:0] R0_data_121_0 = mem_121_0_R0_data;
  wire [7:0] R0_data_121_1 = mem_121_1_R0_data;
  wire [7:0] R0_data_121_2 = mem_121_2_R0_data;
  wire [7:0] R0_data_121_3 = mem_121_3_R0_data;
  wire [7:0] R0_data_121_4 = mem_121_4_R0_data;
  wire [7:0] R0_data_121_5 = mem_121_5_R0_data;
  wire [7:0] R0_data_121_6 = mem_121_6_R0_data;
  wire [7:0] R0_data_121_7 = mem_121_7_R0_data;
  wire [63:0] R0_data_121 = {R0_data_121_7,R0_data_121_6,R0_data_121_5,R0_data_121_4,R0_data_121_3,R0_data_121_2,
    R0_data_121_1,R0_data_121_0};
  wire [7:0] R0_data_122_0 = mem_122_0_R0_data;
  wire [7:0] R0_data_122_1 = mem_122_1_R0_data;
  wire [7:0] R0_data_122_2 = mem_122_2_R0_data;
  wire [7:0] R0_data_122_3 = mem_122_3_R0_data;
  wire [7:0] R0_data_122_4 = mem_122_4_R0_data;
  wire [7:0] R0_data_122_5 = mem_122_5_R0_data;
  wire [7:0] R0_data_122_6 = mem_122_6_R0_data;
  wire [7:0] R0_data_122_7 = mem_122_7_R0_data;
  wire [63:0] R0_data_122 = {R0_data_122_7,R0_data_122_6,R0_data_122_5,R0_data_122_4,R0_data_122_3,R0_data_122_2,
    R0_data_122_1,R0_data_122_0};
  wire [7:0] R0_data_123_0 = mem_123_0_R0_data;
  wire [7:0] R0_data_123_1 = mem_123_1_R0_data;
  wire [7:0] R0_data_123_2 = mem_123_2_R0_data;
  wire [7:0] R0_data_123_3 = mem_123_3_R0_data;
  wire [7:0] R0_data_123_4 = mem_123_4_R0_data;
  wire [7:0] R0_data_123_5 = mem_123_5_R0_data;
  wire [7:0] R0_data_123_6 = mem_123_6_R0_data;
  wire [7:0] R0_data_123_7 = mem_123_7_R0_data;
  wire [63:0] R0_data_123 = {R0_data_123_7,R0_data_123_6,R0_data_123_5,R0_data_123_4,R0_data_123_3,R0_data_123_2,
    R0_data_123_1,R0_data_123_0};
  wire [7:0] R0_data_124_0 = mem_124_0_R0_data;
  wire [7:0] R0_data_124_1 = mem_124_1_R0_data;
  wire [7:0] R0_data_124_2 = mem_124_2_R0_data;
  wire [7:0] R0_data_124_3 = mem_124_3_R0_data;
  wire [7:0] R0_data_124_4 = mem_124_4_R0_data;
  wire [7:0] R0_data_124_5 = mem_124_5_R0_data;
  wire [7:0] R0_data_124_6 = mem_124_6_R0_data;
  wire [7:0] R0_data_124_7 = mem_124_7_R0_data;
  wire [63:0] R0_data_124 = {R0_data_124_7,R0_data_124_6,R0_data_124_5,R0_data_124_4,R0_data_124_3,R0_data_124_2,
    R0_data_124_1,R0_data_124_0};
  wire [7:0] R0_data_125_0 = mem_125_0_R0_data;
  wire [7:0] R0_data_125_1 = mem_125_1_R0_data;
  wire [7:0] R0_data_125_2 = mem_125_2_R0_data;
  wire [7:0] R0_data_125_3 = mem_125_3_R0_data;
  wire [7:0] R0_data_125_4 = mem_125_4_R0_data;
  wire [7:0] R0_data_125_5 = mem_125_5_R0_data;
  wire [7:0] R0_data_125_6 = mem_125_6_R0_data;
  wire [7:0] R0_data_125_7 = mem_125_7_R0_data;
  wire [63:0] R0_data_125 = {R0_data_125_7,R0_data_125_6,R0_data_125_5,R0_data_125_4,R0_data_125_3,R0_data_125_2,
    R0_data_125_1,R0_data_125_0};
  wire [7:0] R0_data_126_0 = mem_126_0_R0_data;
  wire [7:0] R0_data_126_1 = mem_126_1_R0_data;
  wire [7:0] R0_data_126_2 = mem_126_2_R0_data;
  wire [7:0] R0_data_126_3 = mem_126_3_R0_data;
  wire [7:0] R0_data_126_4 = mem_126_4_R0_data;
  wire [7:0] R0_data_126_5 = mem_126_5_R0_data;
  wire [7:0] R0_data_126_6 = mem_126_6_R0_data;
  wire [7:0] R0_data_126_7 = mem_126_7_R0_data;
  wire [63:0] R0_data_126 = {R0_data_126_7,R0_data_126_6,R0_data_126_5,R0_data_126_4,R0_data_126_3,R0_data_126_2,
    R0_data_126_1,R0_data_126_0};
  wire [7:0] R0_data_127_0 = mem_127_0_R0_data;
  wire [7:0] R0_data_127_1 = mem_127_1_R0_data;
  wire [7:0] R0_data_127_2 = mem_127_2_R0_data;
  wire [7:0] R0_data_127_3 = mem_127_3_R0_data;
  wire [7:0] R0_data_127_4 = mem_127_4_R0_data;
  wire [7:0] R0_data_127_5 = mem_127_5_R0_data;
  wire [7:0] R0_data_127_6 = mem_127_6_R0_data;
  wire [7:0] R0_data_127_7 = mem_127_7_R0_data;
  wire [63:0] R0_data_127 = {R0_data_127_7,R0_data_127_6,R0_data_127_5,R0_data_127_4,R0_data_127_3,R0_data_127_2,
    R0_data_127_1,R0_data_127_0};
  wire [7:0] R0_data_128_0 = mem_128_0_R0_data;
  wire [7:0] R0_data_128_1 = mem_128_1_R0_data;
  wire [7:0] R0_data_128_2 = mem_128_2_R0_data;
  wire [7:0] R0_data_128_3 = mem_128_3_R0_data;
  wire [7:0] R0_data_128_4 = mem_128_4_R0_data;
  wire [7:0] R0_data_128_5 = mem_128_5_R0_data;
  wire [7:0] R0_data_128_6 = mem_128_6_R0_data;
  wire [7:0] R0_data_128_7 = mem_128_7_R0_data;
  wire [63:0] R0_data_128 = {R0_data_128_7,R0_data_128_6,R0_data_128_5,R0_data_128_4,R0_data_128_3,R0_data_128_2,
    R0_data_128_1,R0_data_128_0};
  wire [7:0] R0_data_129_0 = mem_129_0_R0_data;
  wire [7:0] R0_data_129_1 = mem_129_1_R0_data;
  wire [7:0] R0_data_129_2 = mem_129_2_R0_data;
  wire [7:0] R0_data_129_3 = mem_129_3_R0_data;
  wire [7:0] R0_data_129_4 = mem_129_4_R0_data;
  wire [7:0] R0_data_129_5 = mem_129_5_R0_data;
  wire [7:0] R0_data_129_6 = mem_129_6_R0_data;
  wire [7:0] R0_data_129_7 = mem_129_7_R0_data;
  wire [63:0] R0_data_129 = {R0_data_129_7,R0_data_129_6,R0_data_129_5,R0_data_129_4,R0_data_129_3,R0_data_129_2,
    R0_data_129_1,R0_data_129_0};
  wire [7:0] R0_data_130_0 = mem_130_0_R0_data;
  wire [7:0] R0_data_130_1 = mem_130_1_R0_data;
  wire [7:0] R0_data_130_2 = mem_130_2_R0_data;
  wire [7:0] R0_data_130_3 = mem_130_3_R0_data;
  wire [7:0] R0_data_130_4 = mem_130_4_R0_data;
  wire [7:0] R0_data_130_5 = mem_130_5_R0_data;
  wire [7:0] R0_data_130_6 = mem_130_6_R0_data;
  wire [7:0] R0_data_130_7 = mem_130_7_R0_data;
  wire [63:0] R0_data_130 = {R0_data_130_7,R0_data_130_6,R0_data_130_5,R0_data_130_4,R0_data_130_3,R0_data_130_2,
    R0_data_130_1,R0_data_130_0};
  wire [7:0] R0_data_131_0 = mem_131_0_R0_data;
  wire [7:0] R0_data_131_1 = mem_131_1_R0_data;
  wire [7:0] R0_data_131_2 = mem_131_2_R0_data;
  wire [7:0] R0_data_131_3 = mem_131_3_R0_data;
  wire [7:0] R0_data_131_4 = mem_131_4_R0_data;
  wire [7:0] R0_data_131_5 = mem_131_5_R0_data;
  wire [7:0] R0_data_131_6 = mem_131_6_R0_data;
  wire [7:0] R0_data_131_7 = mem_131_7_R0_data;
  wire [63:0] R0_data_131 = {R0_data_131_7,R0_data_131_6,R0_data_131_5,R0_data_131_4,R0_data_131_3,R0_data_131_2,
    R0_data_131_1,R0_data_131_0};
  wire [7:0] R0_data_132_0 = mem_132_0_R0_data;
  wire [7:0] R0_data_132_1 = mem_132_1_R0_data;
  wire [7:0] R0_data_132_2 = mem_132_2_R0_data;
  wire [7:0] R0_data_132_3 = mem_132_3_R0_data;
  wire [7:0] R0_data_132_4 = mem_132_4_R0_data;
  wire [7:0] R0_data_132_5 = mem_132_5_R0_data;
  wire [7:0] R0_data_132_6 = mem_132_6_R0_data;
  wire [7:0] R0_data_132_7 = mem_132_7_R0_data;
  wire [63:0] R0_data_132 = {R0_data_132_7,R0_data_132_6,R0_data_132_5,R0_data_132_4,R0_data_132_3,R0_data_132_2,
    R0_data_132_1,R0_data_132_0};
  wire [7:0] R0_data_133_0 = mem_133_0_R0_data;
  wire [7:0] R0_data_133_1 = mem_133_1_R0_data;
  wire [7:0] R0_data_133_2 = mem_133_2_R0_data;
  wire [7:0] R0_data_133_3 = mem_133_3_R0_data;
  wire [7:0] R0_data_133_4 = mem_133_4_R0_data;
  wire [7:0] R0_data_133_5 = mem_133_5_R0_data;
  wire [7:0] R0_data_133_6 = mem_133_6_R0_data;
  wire [7:0] R0_data_133_7 = mem_133_7_R0_data;
  wire [63:0] R0_data_133 = {R0_data_133_7,R0_data_133_6,R0_data_133_5,R0_data_133_4,R0_data_133_3,R0_data_133_2,
    R0_data_133_1,R0_data_133_0};
  wire [7:0] R0_data_134_0 = mem_134_0_R0_data;
  wire [7:0] R0_data_134_1 = mem_134_1_R0_data;
  wire [7:0] R0_data_134_2 = mem_134_2_R0_data;
  wire [7:0] R0_data_134_3 = mem_134_3_R0_data;
  wire [7:0] R0_data_134_4 = mem_134_4_R0_data;
  wire [7:0] R0_data_134_5 = mem_134_5_R0_data;
  wire [7:0] R0_data_134_6 = mem_134_6_R0_data;
  wire [7:0] R0_data_134_7 = mem_134_7_R0_data;
  wire [63:0] R0_data_134 = {R0_data_134_7,R0_data_134_6,R0_data_134_5,R0_data_134_4,R0_data_134_3,R0_data_134_2,
    R0_data_134_1,R0_data_134_0};
  wire [7:0] R0_data_135_0 = mem_135_0_R0_data;
  wire [7:0] R0_data_135_1 = mem_135_1_R0_data;
  wire [7:0] R0_data_135_2 = mem_135_2_R0_data;
  wire [7:0] R0_data_135_3 = mem_135_3_R0_data;
  wire [7:0] R0_data_135_4 = mem_135_4_R0_data;
  wire [7:0] R0_data_135_5 = mem_135_5_R0_data;
  wire [7:0] R0_data_135_6 = mem_135_6_R0_data;
  wire [7:0] R0_data_135_7 = mem_135_7_R0_data;
  wire [63:0] R0_data_135 = {R0_data_135_7,R0_data_135_6,R0_data_135_5,R0_data_135_4,R0_data_135_3,R0_data_135_2,
    R0_data_135_1,R0_data_135_0};
  wire [7:0] R0_data_136_0 = mem_136_0_R0_data;
  wire [7:0] R0_data_136_1 = mem_136_1_R0_data;
  wire [7:0] R0_data_136_2 = mem_136_2_R0_data;
  wire [7:0] R0_data_136_3 = mem_136_3_R0_data;
  wire [7:0] R0_data_136_4 = mem_136_4_R0_data;
  wire [7:0] R0_data_136_5 = mem_136_5_R0_data;
  wire [7:0] R0_data_136_6 = mem_136_6_R0_data;
  wire [7:0] R0_data_136_7 = mem_136_7_R0_data;
  wire [63:0] R0_data_136 = {R0_data_136_7,R0_data_136_6,R0_data_136_5,R0_data_136_4,R0_data_136_3,R0_data_136_2,
    R0_data_136_1,R0_data_136_0};
  wire [7:0] R0_data_137_0 = mem_137_0_R0_data;
  wire [7:0] R0_data_137_1 = mem_137_1_R0_data;
  wire [7:0] R0_data_137_2 = mem_137_2_R0_data;
  wire [7:0] R0_data_137_3 = mem_137_3_R0_data;
  wire [7:0] R0_data_137_4 = mem_137_4_R0_data;
  wire [7:0] R0_data_137_5 = mem_137_5_R0_data;
  wire [7:0] R0_data_137_6 = mem_137_6_R0_data;
  wire [7:0] R0_data_137_7 = mem_137_7_R0_data;
  wire [63:0] R0_data_137 = {R0_data_137_7,R0_data_137_6,R0_data_137_5,R0_data_137_4,R0_data_137_3,R0_data_137_2,
    R0_data_137_1,R0_data_137_0};
  wire [7:0] R0_data_138_0 = mem_138_0_R0_data;
  wire [7:0] R0_data_138_1 = mem_138_1_R0_data;
  wire [7:0] R0_data_138_2 = mem_138_2_R0_data;
  wire [7:0] R0_data_138_3 = mem_138_3_R0_data;
  wire [7:0] R0_data_138_4 = mem_138_4_R0_data;
  wire [7:0] R0_data_138_5 = mem_138_5_R0_data;
  wire [7:0] R0_data_138_6 = mem_138_6_R0_data;
  wire [7:0] R0_data_138_7 = mem_138_7_R0_data;
  wire [63:0] R0_data_138 = {R0_data_138_7,R0_data_138_6,R0_data_138_5,R0_data_138_4,R0_data_138_3,R0_data_138_2,
    R0_data_138_1,R0_data_138_0};
  wire [7:0] R0_data_139_0 = mem_139_0_R0_data;
  wire [7:0] R0_data_139_1 = mem_139_1_R0_data;
  wire [7:0] R0_data_139_2 = mem_139_2_R0_data;
  wire [7:0] R0_data_139_3 = mem_139_3_R0_data;
  wire [7:0] R0_data_139_4 = mem_139_4_R0_data;
  wire [7:0] R0_data_139_5 = mem_139_5_R0_data;
  wire [7:0] R0_data_139_6 = mem_139_6_R0_data;
  wire [7:0] R0_data_139_7 = mem_139_7_R0_data;
  wire [63:0] R0_data_139 = {R0_data_139_7,R0_data_139_6,R0_data_139_5,R0_data_139_4,R0_data_139_3,R0_data_139_2,
    R0_data_139_1,R0_data_139_0};
  wire [7:0] R0_data_140_0 = mem_140_0_R0_data;
  wire [7:0] R0_data_140_1 = mem_140_1_R0_data;
  wire [7:0] R0_data_140_2 = mem_140_2_R0_data;
  wire [7:0] R0_data_140_3 = mem_140_3_R0_data;
  wire [7:0] R0_data_140_4 = mem_140_4_R0_data;
  wire [7:0] R0_data_140_5 = mem_140_5_R0_data;
  wire [7:0] R0_data_140_6 = mem_140_6_R0_data;
  wire [7:0] R0_data_140_7 = mem_140_7_R0_data;
  wire [63:0] R0_data_140 = {R0_data_140_7,R0_data_140_6,R0_data_140_5,R0_data_140_4,R0_data_140_3,R0_data_140_2,
    R0_data_140_1,R0_data_140_0};
  wire [7:0] R0_data_141_0 = mem_141_0_R0_data;
  wire [7:0] R0_data_141_1 = mem_141_1_R0_data;
  wire [7:0] R0_data_141_2 = mem_141_2_R0_data;
  wire [7:0] R0_data_141_3 = mem_141_3_R0_data;
  wire [7:0] R0_data_141_4 = mem_141_4_R0_data;
  wire [7:0] R0_data_141_5 = mem_141_5_R0_data;
  wire [7:0] R0_data_141_6 = mem_141_6_R0_data;
  wire [7:0] R0_data_141_7 = mem_141_7_R0_data;
  wire [63:0] R0_data_141 = {R0_data_141_7,R0_data_141_6,R0_data_141_5,R0_data_141_4,R0_data_141_3,R0_data_141_2,
    R0_data_141_1,R0_data_141_0};
  wire [7:0] R0_data_142_0 = mem_142_0_R0_data;
  wire [7:0] R0_data_142_1 = mem_142_1_R0_data;
  wire [7:0] R0_data_142_2 = mem_142_2_R0_data;
  wire [7:0] R0_data_142_3 = mem_142_3_R0_data;
  wire [7:0] R0_data_142_4 = mem_142_4_R0_data;
  wire [7:0] R0_data_142_5 = mem_142_5_R0_data;
  wire [7:0] R0_data_142_6 = mem_142_6_R0_data;
  wire [7:0] R0_data_142_7 = mem_142_7_R0_data;
  wire [63:0] R0_data_142 = {R0_data_142_7,R0_data_142_6,R0_data_142_5,R0_data_142_4,R0_data_142_3,R0_data_142_2,
    R0_data_142_1,R0_data_142_0};
  wire [7:0] R0_data_143_0 = mem_143_0_R0_data;
  wire [7:0] R0_data_143_1 = mem_143_1_R0_data;
  wire [7:0] R0_data_143_2 = mem_143_2_R0_data;
  wire [7:0] R0_data_143_3 = mem_143_3_R0_data;
  wire [7:0] R0_data_143_4 = mem_143_4_R0_data;
  wire [7:0] R0_data_143_5 = mem_143_5_R0_data;
  wire [7:0] R0_data_143_6 = mem_143_6_R0_data;
  wire [7:0] R0_data_143_7 = mem_143_7_R0_data;
  wire [63:0] R0_data_143 = {R0_data_143_7,R0_data_143_6,R0_data_143_5,R0_data_143_4,R0_data_143_3,R0_data_143_2,
    R0_data_143_1,R0_data_143_0};
  wire [7:0] R0_data_144_0 = mem_144_0_R0_data;
  wire [7:0] R0_data_144_1 = mem_144_1_R0_data;
  wire [7:0] R0_data_144_2 = mem_144_2_R0_data;
  wire [7:0] R0_data_144_3 = mem_144_3_R0_data;
  wire [7:0] R0_data_144_4 = mem_144_4_R0_data;
  wire [7:0] R0_data_144_5 = mem_144_5_R0_data;
  wire [7:0] R0_data_144_6 = mem_144_6_R0_data;
  wire [7:0] R0_data_144_7 = mem_144_7_R0_data;
  wire [63:0] R0_data_144 = {R0_data_144_7,R0_data_144_6,R0_data_144_5,R0_data_144_4,R0_data_144_3,R0_data_144_2,
    R0_data_144_1,R0_data_144_0};
  wire [7:0] R0_data_145_0 = mem_145_0_R0_data;
  wire [7:0] R0_data_145_1 = mem_145_1_R0_data;
  wire [7:0] R0_data_145_2 = mem_145_2_R0_data;
  wire [7:0] R0_data_145_3 = mem_145_3_R0_data;
  wire [7:0] R0_data_145_4 = mem_145_4_R0_data;
  wire [7:0] R0_data_145_5 = mem_145_5_R0_data;
  wire [7:0] R0_data_145_6 = mem_145_6_R0_data;
  wire [7:0] R0_data_145_7 = mem_145_7_R0_data;
  wire [63:0] R0_data_145 = {R0_data_145_7,R0_data_145_6,R0_data_145_5,R0_data_145_4,R0_data_145_3,R0_data_145_2,
    R0_data_145_1,R0_data_145_0};
  wire [7:0] R0_data_146_0 = mem_146_0_R0_data;
  wire [7:0] R0_data_146_1 = mem_146_1_R0_data;
  wire [7:0] R0_data_146_2 = mem_146_2_R0_data;
  wire [7:0] R0_data_146_3 = mem_146_3_R0_data;
  wire [7:0] R0_data_146_4 = mem_146_4_R0_data;
  wire [7:0] R0_data_146_5 = mem_146_5_R0_data;
  wire [7:0] R0_data_146_6 = mem_146_6_R0_data;
  wire [7:0] R0_data_146_7 = mem_146_7_R0_data;
  wire [63:0] R0_data_146 = {R0_data_146_7,R0_data_146_6,R0_data_146_5,R0_data_146_4,R0_data_146_3,R0_data_146_2,
    R0_data_146_1,R0_data_146_0};
  wire [7:0] R0_data_147_0 = mem_147_0_R0_data;
  wire [7:0] R0_data_147_1 = mem_147_1_R0_data;
  wire [7:0] R0_data_147_2 = mem_147_2_R0_data;
  wire [7:0] R0_data_147_3 = mem_147_3_R0_data;
  wire [7:0] R0_data_147_4 = mem_147_4_R0_data;
  wire [7:0] R0_data_147_5 = mem_147_5_R0_data;
  wire [7:0] R0_data_147_6 = mem_147_6_R0_data;
  wire [7:0] R0_data_147_7 = mem_147_7_R0_data;
  wire [63:0] R0_data_147 = {R0_data_147_7,R0_data_147_6,R0_data_147_5,R0_data_147_4,R0_data_147_3,R0_data_147_2,
    R0_data_147_1,R0_data_147_0};
  wire [7:0] R0_data_148_0 = mem_148_0_R0_data;
  wire [7:0] R0_data_148_1 = mem_148_1_R0_data;
  wire [7:0] R0_data_148_2 = mem_148_2_R0_data;
  wire [7:0] R0_data_148_3 = mem_148_3_R0_data;
  wire [7:0] R0_data_148_4 = mem_148_4_R0_data;
  wire [7:0] R0_data_148_5 = mem_148_5_R0_data;
  wire [7:0] R0_data_148_6 = mem_148_6_R0_data;
  wire [7:0] R0_data_148_7 = mem_148_7_R0_data;
  wire [63:0] R0_data_148 = {R0_data_148_7,R0_data_148_6,R0_data_148_5,R0_data_148_4,R0_data_148_3,R0_data_148_2,
    R0_data_148_1,R0_data_148_0};
  wire [7:0] R0_data_149_0 = mem_149_0_R0_data;
  wire [7:0] R0_data_149_1 = mem_149_1_R0_data;
  wire [7:0] R0_data_149_2 = mem_149_2_R0_data;
  wire [7:0] R0_data_149_3 = mem_149_3_R0_data;
  wire [7:0] R0_data_149_4 = mem_149_4_R0_data;
  wire [7:0] R0_data_149_5 = mem_149_5_R0_data;
  wire [7:0] R0_data_149_6 = mem_149_6_R0_data;
  wire [7:0] R0_data_149_7 = mem_149_7_R0_data;
  wire [63:0] R0_data_149 = {R0_data_149_7,R0_data_149_6,R0_data_149_5,R0_data_149_4,R0_data_149_3,R0_data_149_2,
    R0_data_149_1,R0_data_149_0};
  wire [7:0] R0_data_150_0 = mem_150_0_R0_data;
  wire [7:0] R0_data_150_1 = mem_150_1_R0_data;
  wire [7:0] R0_data_150_2 = mem_150_2_R0_data;
  wire [7:0] R0_data_150_3 = mem_150_3_R0_data;
  wire [7:0] R0_data_150_4 = mem_150_4_R0_data;
  wire [7:0] R0_data_150_5 = mem_150_5_R0_data;
  wire [7:0] R0_data_150_6 = mem_150_6_R0_data;
  wire [7:0] R0_data_150_7 = mem_150_7_R0_data;
  wire [63:0] R0_data_150 = {R0_data_150_7,R0_data_150_6,R0_data_150_5,R0_data_150_4,R0_data_150_3,R0_data_150_2,
    R0_data_150_1,R0_data_150_0};
  wire [7:0] R0_data_151_0 = mem_151_0_R0_data;
  wire [7:0] R0_data_151_1 = mem_151_1_R0_data;
  wire [7:0] R0_data_151_2 = mem_151_2_R0_data;
  wire [7:0] R0_data_151_3 = mem_151_3_R0_data;
  wire [7:0] R0_data_151_4 = mem_151_4_R0_data;
  wire [7:0] R0_data_151_5 = mem_151_5_R0_data;
  wire [7:0] R0_data_151_6 = mem_151_6_R0_data;
  wire [7:0] R0_data_151_7 = mem_151_7_R0_data;
  wire [63:0] R0_data_151 = {R0_data_151_7,R0_data_151_6,R0_data_151_5,R0_data_151_4,R0_data_151_3,R0_data_151_2,
    R0_data_151_1,R0_data_151_0};
  wire [7:0] R0_data_152_0 = mem_152_0_R0_data;
  wire [7:0] R0_data_152_1 = mem_152_1_R0_data;
  wire [7:0] R0_data_152_2 = mem_152_2_R0_data;
  wire [7:0] R0_data_152_3 = mem_152_3_R0_data;
  wire [7:0] R0_data_152_4 = mem_152_4_R0_data;
  wire [7:0] R0_data_152_5 = mem_152_5_R0_data;
  wire [7:0] R0_data_152_6 = mem_152_6_R0_data;
  wire [7:0] R0_data_152_7 = mem_152_7_R0_data;
  wire [63:0] R0_data_152 = {R0_data_152_7,R0_data_152_6,R0_data_152_5,R0_data_152_4,R0_data_152_3,R0_data_152_2,
    R0_data_152_1,R0_data_152_0};
  wire [7:0] R0_data_153_0 = mem_153_0_R0_data;
  wire [7:0] R0_data_153_1 = mem_153_1_R0_data;
  wire [7:0] R0_data_153_2 = mem_153_2_R0_data;
  wire [7:0] R0_data_153_3 = mem_153_3_R0_data;
  wire [7:0] R0_data_153_4 = mem_153_4_R0_data;
  wire [7:0] R0_data_153_5 = mem_153_5_R0_data;
  wire [7:0] R0_data_153_6 = mem_153_6_R0_data;
  wire [7:0] R0_data_153_7 = mem_153_7_R0_data;
  wire [63:0] R0_data_153 = {R0_data_153_7,R0_data_153_6,R0_data_153_5,R0_data_153_4,R0_data_153_3,R0_data_153_2,
    R0_data_153_1,R0_data_153_0};
  wire [7:0] R0_data_154_0 = mem_154_0_R0_data;
  wire [7:0] R0_data_154_1 = mem_154_1_R0_data;
  wire [7:0] R0_data_154_2 = mem_154_2_R0_data;
  wire [7:0] R0_data_154_3 = mem_154_3_R0_data;
  wire [7:0] R0_data_154_4 = mem_154_4_R0_data;
  wire [7:0] R0_data_154_5 = mem_154_5_R0_data;
  wire [7:0] R0_data_154_6 = mem_154_6_R0_data;
  wire [7:0] R0_data_154_7 = mem_154_7_R0_data;
  wire [63:0] R0_data_154 = {R0_data_154_7,R0_data_154_6,R0_data_154_5,R0_data_154_4,R0_data_154_3,R0_data_154_2,
    R0_data_154_1,R0_data_154_0};
  wire [7:0] R0_data_155_0 = mem_155_0_R0_data;
  wire [7:0] R0_data_155_1 = mem_155_1_R0_data;
  wire [7:0] R0_data_155_2 = mem_155_2_R0_data;
  wire [7:0] R0_data_155_3 = mem_155_3_R0_data;
  wire [7:0] R0_data_155_4 = mem_155_4_R0_data;
  wire [7:0] R0_data_155_5 = mem_155_5_R0_data;
  wire [7:0] R0_data_155_6 = mem_155_6_R0_data;
  wire [7:0] R0_data_155_7 = mem_155_7_R0_data;
  wire [63:0] R0_data_155 = {R0_data_155_7,R0_data_155_6,R0_data_155_5,R0_data_155_4,R0_data_155_3,R0_data_155_2,
    R0_data_155_1,R0_data_155_0};
  wire [7:0] R0_data_156_0 = mem_156_0_R0_data;
  wire [7:0] R0_data_156_1 = mem_156_1_R0_data;
  wire [7:0] R0_data_156_2 = mem_156_2_R0_data;
  wire [7:0] R0_data_156_3 = mem_156_3_R0_data;
  wire [7:0] R0_data_156_4 = mem_156_4_R0_data;
  wire [7:0] R0_data_156_5 = mem_156_5_R0_data;
  wire [7:0] R0_data_156_6 = mem_156_6_R0_data;
  wire [7:0] R0_data_156_7 = mem_156_7_R0_data;
  wire [63:0] R0_data_156 = {R0_data_156_7,R0_data_156_6,R0_data_156_5,R0_data_156_4,R0_data_156_3,R0_data_156_2,
    R0_data_156_1,R0_data_156_0};
  wire [7:0] R0_data_157_0 = mem_157_0_R0_data;
  wire [7:0] R0_data_157_1 = mem_157_1_R0_data;
  wire [7:0] R0_data_157_2 = mem_157_2_R0_data;
  wire [7:0] R0_data_157_3 = mem_157_3_R0_data;
  wire [7:0] R0_data_157_4 = mem_157_4_R0_data;
  wire [7:0] R0_data_157_5 = mem_157_5_R0_data;
  wire [7:0] R0_data_157_6 = mem_157_6_R0_data;
  wire [7:0] R0_data_157_7 = mem_157_7_R0_data;
  wire [63:0] R0_data_157 = {R0_data_157_7,R0_data_157_6,R0_data_157_5,R0_data_157_4,R0_data_157_3,R0_data_157_2,
    R0_data_157_1,R0_data_157_0};
  wire [7:0] R0_data_158_0 = mem_158_0_R0_data;
  wire [7:0] R0_data_158_1 = mem_158_1_R0_data;
  wire [7:0] R0_data_158_2 = mem_158_2_R0_data;
  wire [7:0] R0_data_158_3 = mem_158_3_R0_data;
  wire [7:0] R0_data_158_4 = mem_158_4_R0_data;
  wire [7:0] R0_data_158_5 = mem_158_5_R0_data;
  wire [7:0] R0_data_158_6 = mem_158_6_R0_data;
  wire [7:0] R0_data_158_7 = mem_158_7_R0_data;
  wire [63:0] R0_data_158 = {R0_data_158_7,R0_data_158_6,R0_data_158_5,R0_data_158_4,R0_data_158_3,R0_data_158_2,
    R0_data_158_1,R0_data_158_0};
  wire [7:0] R0_data_159_0 = mem_159_0_R0_data;
  wire [7:0] R0_data_159_1 = mem_159_1_R0_data;
  wire [7:0] R0_data_159_2 = mem_159_2_R0_data;
  wire [7:0] R0_data_159_3 = mem_159_3_R0_data;
  wire [7:0] R0_data_159_4 = mem_159_4_R0_data;
  wire [7:0] R0_data_159_5 = mem_159_5_R0_data;
  wire [7:0] R0_data_159_6 = mem_159_6_R0_data;
  wire [7:0] R0_data_159_7 = mem_159_7_R0_data;
  wire [63:0] R0_data_159 = {R0_data_159_7,R0_data_159_6,R0_data_159_5,R0_data_159_4,R0_data_159_3,R0_data_159_2,
    R0_data_159_1,R0_data_159_0};
  wire [7:0] R0_data_160_0 = mem_160_0_R0_data;
  wire [7:0] R0_data_160_1 = mem_160_1_R0_data;
  wire [7:0] R0_data_160_2 = mem_160_2_R0_data;
  wire [7:0] R0_data_160_3 = mem_160_3_R0_data;
  wire [7:0] R0_data_160_4 = mem_160_4_R0_data;
  wire [7:0] R0_data_160_5 = mem_160_5_R0_data;
  wire [7:0] R0_data_160_6 = mem_160_6_R0_data;
  wire [7:0] R0_data_160_7 = mem_160_7_R0_data;
  wire [63:0] R0_data_160 = {R0_data_160_7,R0_data_160_6,R0_data_160_5,R0_data_160_4,R0_data_160_3,R0_data_160_2,
    R0_data_160_1,R0_data_160_0};
  wire [7:0] R0_data_161_0 = mem_161_0_R0_data;
  wire [7:0] R0_data_161_1 = mem_161_1_R0_data;
  wire [7:0] R0_data_161_2 = mem_161_2_R0_data;
  wire [7:0] R0_data_161_3 = mem_161_3_R0_data;
  wire [7:0] R0_data_161_4 = mem_161_4_R0_data;
  wire [7:0] R0_data_161_5 = mem_161_5_R0_data;
  wire [7:0] R0_data_161_6 = mem_161_6_R0_data;
  wire [7:0] R0_data_161_7 = mem_161_7_R0_data;
  wire [63:0] R0_data_161 = {R0_data_161_7,R0_data_161_6,R0_data_161_5,R0_data_161_4,R0_data_161_3,R0_data_161_2,
    R0_data_161_1,R0_data_161_0};
  wire [7:0] R0_data_162_0 = mem_162_0_R0_data;
  wire [7:0] R0_data_162_1 = mem_162_1_R0_data;
  wire [7:0] R0_data_162_2 = mem_162_2_R0_data;
  wire [7:0] R0_data_162_3 = mem_162_3_R0_data;
  wire [7:0] R0_data_162_4 = mem_162_4_R0_data;
  wire [7:0] R0_data_162_5 = mem_162_5_R0_data;
  wire [7:0] R0_data_162_6 = mem_162_6_R0_data;
  wire [7:0] R0_data_162_7 = mem_162_7_R0_data;
  wire [63:0] R0_data_162 = {R0_data_162_7,R0_data_162_6,R0_data_162_5,R0_data_162_4,R0_data_162_3,R0_data_162_2,
    R0_data_162_1,R0_data_162_0};
  wire [7:0] R0_data_163_0 = mem_163_0_R0_data;
  wire [7:0] R0_data_163_1 = mem_163_1_R0_data;
  wire [7:0] R0_data_163_2 = mem_163_2_R0_data;
  wire [7:0] R0_data_163_3 = mem_163_3_R0_data;
  wire [7:0] R0_data_163_4 = mem_163_4_R0_data;
  wire [7:0] R0_data_163_5 = mem_163_5_R0_data;
  wire [7:0] R0_data_163_6 = mem_163_6_R0_data;
  wire [7:0] R0_data_163_7 = mem_163_7_R0_data;
  wire [63:0] R0_data_163 = {R0_data_163_7,R0_data_163_6,R0_data_163_5,R0_data_163_4,R0_data_163_3,R0_data_163_2,
    R0_data_163_1,R0_data_163_0};
  wire [7:0] R0_data_164_0 = mem_164_0_R0_data;
  wire [7:0] R0_data_164_1 = mem_164_1_R0_data;
  wire [7:0] R0_data_164_2 = mem_164_2_R0_data;
  wire [7:0] R0_data_164_3 = mem_164_3_R0_data;
  wire [7:0] R0_data_164_4 = mem_164_4_R0_data;
  wire [7:0] R0_data_164_5 = mem_164_5_R0_data;
  wire [7:0] R0_data_164_6 = mem_164_6_R0_data;
  wire [7:0] R0_data_164_7 = mem_164_7_R0_data;
  wire [63:0] R0_data_164 = {R0_data_164_7,R0_data_164_6,R0_data_164_5,R0_data_164_4,R0_data_164_3,R0_data_164_2,
    R0_data_164_1,R0_data_164_0};
  wire [7:0] R0_data_165_0 = mem_165_0_R0_data;
  wire [7:0] R0_data_165_1 = mem_165_1_R0_data;
  wire [7:0] R0_data_165_2 = mem_165_2_R0_data;
  wire [7:0] R0_data_165_3 = mem_165_3_R0_data;
  wire [7:0] R0_data_165_4 = mem_165_4_R0_data;
  wire [7:0] R0_data_165_5 = mem_165_5_R0_data;
  wire [7:0] R0_data_165_6 = mem_165_6_R0_data;
  wire [7:0] R0_data_165_7 = mem_165_7_R0_data;
  wire [63:0] R0_data_165 = {R0_data_165_7,R0_data_165_6,R0_data_165_5,R0_data_165_4,R0_data_165_3,R0_data_165_2,
    R0_data_165_1,R0_data_165_0};
  wire [7:0] R0_data_166_0 = mem_166_0_R0_data;
  wire [7:0] R0_data_166_1 = mem_166_1_R0_data;
  wire [7:0] R0_data_166_2 = mem_166_2_R0_data;
  wire [7:0] R0_data_166_3 = mem_166_3_R0_data;
  wire [7:0] R0_data_166_4 = mem_166_4_R0_data;
  wire [7:0] R0_data_166_5 = mem_166_5_R0_data;
  wire [7:0] R0_data_166_6 = mem_166_6_R0_data;
  wire [7:0] R0_data_166_7 = mem_166_7_R0_data;
  wire [63:0] R0_data_166 = {R0_data_166_7,R0_data_166_6,R0_data_166_5,R0_data_166_4,R0_data_166_3,R0_data_166_2,
    R0_data_166_1,R0_data_166_0};
  wire [7:0] R0_data_167_0 = mem_167_0_R0_data;
  wire [7:0] R0_data_167_1 = mem_167_1_R0_data;
  wire [7:0] R0_data_167_2 = mem_167_2_R0_data;
  wire [7:0] R0_data_167_3 = mem_167_3_R0_data;
  wire [7:0] R0_data_167_4 = mem_167_4_R0_data;
  wire [7:0] R0_data_167_5 = mem_167_5_R0_data;
  wire [7:0] R0_data_167_6 = mem_167_6_R0_data;
  wire [7:0] R0_data_167_7 = mem_167_7_R0_data;
  wire [63:0] R0_data_167 = {R0_data_167_7,R0_data_167_6,R0_data_167_5,R0_data_167_4,R0_data_167_3,R0_data_167_2,
    R0_data_167_1,R0_data_167_0};
  wire [7:0] R0_data_168_0 = mem_168_0_R0_data;
  wire [7:0] R0_data_168_1 = mem_168_1_R0_data;
  wire [7:0] R0_data_168_2 = mem_168_2_R0_data;
  wire [7:0] R0_data_168_3 = mem_168_3_R0_data;
  wire [7:0] R0_data_168_4 = mem_168_4_R0_data;
  wire [7:0] R0_data_168_5 = mem_168_5_R0_data;
  wire [7:0] R0_data_168_6 = mem_168_6_R0_data;
  wire [7:0] R0_data_168_7 = mem_168_7_R0_data;
  wire [63:0] R0_data_168 = {R0_data_168_7,R0_data_168_6,R0_data_168_5,R0_data_168_4,R0_data_168_3,R0_data_168_2,
    R0_data_168_1,R0_data_168_0};
  wire [7:0] R0_data_169_0 = mem_169_0_R0_data;
  wire [7:0] R0_data_169_1 = mem_169_1_R0_data;
  wire [7:0] R0_data_169_2 = mem_169_2_R0_data;
  wire [7:0] R0_data_169_3 = mem_169_3_R0_data;
  wire [7:0] R0_data_169_4 = mem_169_4_R0_data;
  wire [7:0] R0_data_169_5 = mem_169_5_R0_data;
  wire [7:0] R0_data_169_6 = mem_169_6_R0_data;
  wire [7:0] R0_data_169_7 = mem_169_7_R0_data;
  wire [63:0] R0_data_169 = {R0_data_169_7,R0_data_169_6,R0_data_169_5,R0_data_169_4,R0_data_169_3,R0_data_169_2,
    R0_data_169_1,R0_data_169_0};
  wire [7:0] R0_data_170_0 = mem_170_0_R0_data;
  wire [7:0] R0_data_170_1 = mem_170_1_R0_data;
  wire [7:0] R0_data_170_2 = mem_170_2_R0_data;
  wire [7:0] R0_data_170_3 = mem_170_3_R0_data;
  wire [7:0] R0_data_170_4 = mem_170_4_R0_data;
  wire [7:0] R0_data_170_5 = mem_170_5_R0_data;
  wire [7:0] R0_data_170_6 = mem_170_6_R0_data;
  wire [7:0] R0_data_170_7 = mem_170_7_R0_data;
  wire [63:0] R0_data_170 = {R0_data_170_7,R0_data_170_6,R0_data_170_5,R0_data_170_4,R0_data_170_3,R0_data_170_2,
    R0_data_170_1,R0_data_170_0};
  wire [7:0] R0_data_171_0 = mem_171_0_R0_data;
  wire [7:0] R0_data_171_1 = mem_171_1_R0_data;
  wire [7:0] R0_data_171_2 = mem_171_2_R0_data;
  wire [7:0] R0_data_171_3 = mem_171_3_R0_data;
  wire [7:0] R0_data_171_4 = mem_171_4_R0_data;
  wire [7:0] R0_data_171_5 = mem_171_5_R0_data;
  wire [7:0] R0_data_171_6 = mem_171_6_R0_data;
  wire [7:0] R0_data_171_7 = mem_171_7_R0_data;
  wire [63:0] R0_data_171 = {R0_data_171_7,R0_data_171_6,R0_data_171_5,R0_data_171_4,R0_data_171_3,R0_data_171_2,
    R0_data_171_1,R0_data_171_0};
  wire [7:0] R0_data_172_0 = mem_172_0_R0_data;
  wire [7:0] R0_data_172_1 = mem_172_1_R0_data;
  wire [7:0] R0_data_172_2 = mem_172_2_R0_data;
  wire [7:0] R0_data_172_3 = mem_172_3_R0_data;
  wire [7:0] R0_data_172_4 = mem_172_4_R0_data;
  wire [7:0] R0_data_172_5 = mem_172_5_R0_data;
  wire [7:0] R0_data_172_6 = mem_172_6_R0_data;
  wire [7:0] R0_data_172_7 = mem_172_7_R0_data;
  wire [63:0] R0_data_172 = {R0_data_172_7,R0_data_172_6,R0_data_172_5,R0_data_172_4,R0_data_172_3,R0_data_172_2,
    R0_data_172_1,R0_data_172_0};
  wire [7:0] R0_data_173_0 = mem_173_0_R0_data;
  wire [7:0] R0_data_173_1 = mem_173_1_R0_data;
  wire [7:0] R0_data_173_2 = mem_173_2_R0_data;
  wire [7:0] R0_data_173_3 = mem_173_3_R0_data;
  wire [7:0] R0_data_173_4 = mem_173_4_R0_data;
  wire [7:0] R0_data_173_5 = mem_173_5_R0_data;
  wire [7:0] R0_data_173_6 = mem_173_6_R0_data;
  wire [7:0] R0_data_173_7 = mem_173_7_R0_data;
  wire [63:0] R0_data_173 = {R0_data_173_7,R0_data_173_6,R0_data_173_5,R0_data_173_4,R0_data_173_3,R0_data_173_2,
    R0_data_173_1,R0_data_173_0};
  wire [7:0] R0_data_174_0 = mem_174_0_R0_data;
  wire [7:0] R0_data_174_1 = mem_174_1_R0_data;
  wire [7:0] R0_data_174_2 = mem_174_2_R0_data;
  wire [7:0] R0_data_174_3 = mem_174_3_R0_data;
  wire [7:0] R0_data_174_4 = mem_174_4_R0_data;
  wire [7:0] R0_data_174_5 = mem_174_5_R0_data;
  wire [7:0] R0_data_174_6 = mem_174_6_R0_data;
  wire [7:0] R0_data_174_7 = mem_174_7_R0_data;
  wire [63:0] R0_data_174 = {R0_data_174_7,R0_data_174_6,R0_data_174_5,R0_data_174_4,R0_data_174_3,R0_data_174_2,
    R0_data_174_1,R0_data_174_0};
  wire [7:0] R0_data_175_0 = mem_175_0_R0_data;
  wire [7:0] R0_data_175_1 = mem_175_1_R0_data;
  wire [7:0] R0_data_175_2 = mem_175_2_R0_data;
  wire [7:0] R0_data_175_3 = mem_175_3_R0_data;
  wire [7:0] R0_data_175_4 = mem_175_4_R0_data;
  wire [7:0] R0_data_175_5 = mem_175_5_R0_data;
  wire [7:0] R0_data_175_6 = mem_175_6_R0_data;
  wire [7:0] R0_data_175_7 = mem_175_7_R0_data;
  wire [63:0] R0_data_175 = {R0_data_175_7,R0_data_175_6,R0_data_175_5,R0_data_175_4,R0_data_175_3,R0_data_175_2,
    R0_data_175_1,R0_data_175_0};
  wire [7:0] R0_data_176_0 = mem_176_0_R0_data;
  wire [7:0] R0_data_176_1 = mem_176_1_R0_data;
  wire [7:0] R0_data_176_2 = mem_176_2_R0_data;
  wire [7:0] R0_data_176_3 = mem_176_3_R0_data;
  wire [7:0] R0_data_176_4 = mem_176_4_R0_data;
  wire [7:0] R0_data_176_5 = mem_176_5_R0_data;
  wire [7:0] R0_data_176_6 = mem_176_6_R0_data;
  wire [7:0] R0_data_176_7 = mem_176_7_R0_data;
  wire [63:0] R0_data_176 = {R0_data_176_7,R0_data_176_6,R0_data_176_5,R0_data_176_4,R0_data_176_3,R0_data_176_2,
    R0_data_176_1,R0_data_176_0};
  wire [7:0] R0_data_177_0 = mem_177_0_R0_data;
  wire [7:0] R0_data_177_1 = mem_177_1_R0_data;
  wire [7:0] R0_data_177_2 = mem_177_2_R0_data;
  wire [7:0] R0_data_177_3 = mem_177_3_R0_data;
  wire [7:0] R0_data_177_4 = mem_177_4_R0_data;
  wire [7:0] R0_data_177_5 = mem_177_5_R0_data;
  wire [7:0] R0_data_177_6 = mem_177_6_R0_data;
  wire [7:0] R0_data_177_7 = mem_177_7_R0_data;
  wire [63:0] R0_data_177 = {R0_data_177_7,R0_data_177_6,R0_data_177_5,R0_data_177_4,R0_data_177_3,R0_data_177_2,
    R0_data_177_1,R0_data_177_0};
  wire [7:0] R0_data_178_0 = mem_178_0_R0_data;
  wire [7:0] R0_data_178_1 = mem_178_1_R0_data;
  wire [7:0] R0_data_178_2 = mem_178_2_R0_data;
  wire [7:0] R0_data_178_3 = mem_178_3_R0_data;
  wire [7:0] R0_data_178_4 = mem_178_4_R0_data;
  wire [7:0] R0_data_178_5 = mem_178_5_R0_data;
  wire [7:0] R0_data_178_6 = mem_178_6_R0_data;
  wire [7:0] R0_data_178_7 = mem_178_7_R0_data;
  wire [63:0] R0_data_178 = {R0_data_178_7,R0_data_178_6,R0_data_178_5,R0_data_178_4,R0_data_178_3,R0_data_178_2,
    R0_data_178_1,R0_data_178_0};
  wire [7:0] R0_data_179_0 = mem_179_0_R0_data;
  wire [7:0] R0_data_179_1 = mem_179_1_R0_data;
  wire [7:0] R0_data_179_2 = mem_179_2_R0_data;
  wire [7:0] R0_data_179_3 = mem_179_3_R0_data;
  wire [7:0] R0_data_179_4 = mem_179_4_R0_data;
  wire [7:0] R0_data_179_5 = mem_179_5_R0_data;
  wire [7:0] R0_data_179_6 = mem_179_6_R0_data;
  wire [7:0] R0_data_179_7 = mem_179_7_R0_data;
  wire [63:0] R0_data_179 = {R0_data_179_7,R0_data_179_6,R0_data_179_5,R0_data_179_4,R0_data_179_3,R0_data_179_2,
    R0_data_179_1,R0_data_179_0};
  wire [7:0] R0_data_180_0 = mem_180_0_R0_data;
  wire [7:0] R0_data_180_1 = mem_180_1_R0_data;
  wire [7:0] R0_data_180_2 = mem_180_2_R0_data;
  wire [7:0] R0_data_180_3 = mem_180_3_R0_data;
  wire [7:0] R0_data_180_4 = mem_180_4_R0_data;
  wire [7:0] R0_data_180_5 = mem_180_5_R0_data;
  wire [7:0] R0_data_180_6 = mem_180_6_R0_data;
  wire [7:0] R0_data_180_7 = mem_180_7_R0_data;
  wire [63:0] R0_data_180 = {R0_data_180_7,R0_data_180_6,R0_data_180_5,R0_data_180_4,R0_data_180_3,R0_data_180_2,
    R0_data_180_1,R0_data_180_0};
  wire [7:0] R0_data_181_0 = mem_181_0_R0_data;
  wire [7:0] R0_data_181_1 = mem_181_1_R0_data;
  wire [7:0] R0_data_181_2 = mem_181_2_R0_data;
  wire [7:0] R0_data_181_3 = mem_181_3_R0_data;
  wire [7:0] R0_data_181_4 = mem_181_4_R0_data;
  wire [7:0] R0_data_181_5 = mem_181_5_R0_data;
  wire [7:0] R0_data_181_6 = mem_181_6_R0_data;
  wire [7:0] R0_data_181_7 = mem_181_7_R0_data;
  wire [63:0] R0_data_181 = {R0_data_181_7,R0_data_181_6,R0_data_181_5,R0_data_181_4,R0_data_181_3,R0_data_181_2,
    R0_data_181_1,R0_data_181_0};
  wire [7:0] R0_data_182_0 = mem_182_0_R0_data;
  wire [7:0] R0_data_182_1 = mem_182_1_R0_data;
  wire [7:0] R0_data_182_2 = mem_182_2_R0_data;
  wire [7:0] R0_data_182_3 = mem_182_3_R0_data;
  wire [7:0] R0_data_182_4 = mem_182_4_R0_data;
  wire [7:0] R0_data_182_5 = mem_182_5_R0_data;
  wire [7:0] R0_data_182_6 = mem_182_6_R0_data;
  wire [7:0] R0_data_182_7 = mem_182_7_R0_data;
  wire [63:0] R0_data_182 = {R0_data_182_7,R0_data_182_6,R0_data_182_5,R0_data_182_4,R0_data_182_3,R0_data_182_2,
    R0_data_182_1,R0_data_182_0};
  wire [7:0] R0_data_183_0 = mem_183_0_R0_data;
  wire [7:0] R0_data_183_1 = mem_183_1_R0_data;
  wire [7:0] R0_data_183_2 = mem_183_2_R0_data;
  wire [7:0] R0_data_183_3 = mem_183_3_R0_data;
  wire [7:0] R0_data_183_4 = mem_183_4_R0_data;
  wire [7:0] R0_data_183_5 = mem_183_5_R0_data;
  wire [7:0] R0_data_183_6 = mem_183_6_R0_data;
  wire [7:0] R0_data_183_7 = mem_183_7_R0_data;
  wire [63:0] R0_data_183 = {R0_data_183_7,R0_data_183_6,R0_data_183_5,R0_data_183_4,R0_data_183_3,R0_data_183_2,
    R0_data_183_1,R0_data_183_0};
  wire [7:0] R0_data_184_0 = mem_184_0_R0_data;
  wire [7:0] R0_data_184_1 = mem_184_1_R0_data;
  wire [7:0] R0_data_184_2 = mem_184_2_R0_data;
  wire [7:0] R0_data_184_3 = mem_184_3_R0_data;
  wire [7:0] R0_data_184_4 = mem_184_4_R0_data;
  wire [7:0] R0_data_184_5 = mem_184_5_R0_data;
  wire [7:0] R0_data_184_6 = mem_184_6_R0_data;
  wire [7:0] R0_data_184_7 = mem_184_7_R0_data;
  wire [63:0] R0_data_184 = {R0_data_184_7,R0_data_184_6,R0_data_184_5,R0_data_184_4,R0_data_184_3,R0_data_184_2,
    R0_data_184_1,R0_data_184_0};
  wire [7:0] R0_data_185_0 = mem_185_0_R0_data;
  wire [7:0] R0_data_185_1 = mem_185_1_R0_data;
  wire [7:0] R0_data_185_2 = mem_185_2_R0_data;
  wire [7:0] R0_data_185_3 = mem_185_3_R0_data;
  wire [7:0] R0_data_185_4 = mem_185_4_R0_data;
  wire [7:0] R0_data_185_5 = mem_185_5_R0_data;
  wire [7:0] R0_data_185_6 = mem_185_6_R0_data;
  wire [7:0] R0_data_185_7 = mem_185_7_R0_data;
  wire [63:0] R0_data_185 = {R0_data_185_7,R0_data_185_6,R0_data_185_5,R0_data_185_4,R0_data_185_3,R0_data_185_2,
    R0_data_185_1,R0_data_185_0};
  wire [7:0] R0_data_186_0 = mem_186_0_R0_data;
  wire [7:0] R0_data_186_1 = mem_186_1_R0_data;
  wire [7:0] R0_data_186_2 = mem_186_2_R0_data;
  wire [7:0] R0_data_186_3 = mem_186_3_R0_data;
  wire [7:0] R0_data_186_4 = mem_186_4_R0_data;
  wire [7:0] R0_data_186_5 = mem_186_5_R0_data;
  wire [7:0] R0_data_186_6 = mem_186_6_R0_data;
  wire [7:0] R0_data_186_7 = mem_186_7_R0_data;
  wire [63:0] R0_data_186 = {R0_data_186_7,R0_data_186_6,R0_data_186_5,R0_data_186_4,R0_data_186_3,R0_data_186_2,
    R0_data_186_1,R0_data_186_0};
  wire [7:0] R0_data_187_0 = mem_187_0_R0_data;
  wire [7:0] R0_data_187_1 = mem_187_1_R0_data;
  wire [7:0] R0_data_187_2 = mem_187_2_R0_data;
  wire [7:0] R0_data_187_3 = mem_187_3_R0_data;
  wire [7:0] R0_data_187_4 = mem_187_4_R0_data;
  wire [7:0] R0_data_187_5 = mem_187_5_R0_data;
  wire [7:0] R0_data_187_6 = mem_187_6_R0_data;
  wire [7:0] R0_data_187_7 = mem_187_7_R0_data;
  wire [63:0] R0_data_187 = {R0_data_187_7,R0_data_187_6,R0_data_187_5,R0_data_187_4,R0_data_187_3,R0_data_187_2,
    R0_data_187_1,R0_data_187_0};
  wire [7:0] R0_data_188_0 = mem_188_0_R0_data;
  wire [7:0] R0_data_188_1 = mem_188_1_R0_data;
  wire [7:0] R0_data_188_2 = mem_188_2_R0_data;
  wire [7:0] R0_data_188_3 = mem_188_3_R0_data;
  wire [7:0] R0_data_188_4 = mem_188_4_R0_data;
  wire [7:0] R0_data_188_5 = mem_188_5_R0_data;
  wire [7:0] R0_data_188_6 = mem_188_6_R0_data;
  wire [7:0] R0_data_188_7 = mem_188_7_R0_data;
  wire [63:0] R0_data_188 = {R0_data_188_7,R0_data_188_6,R0_data_188_5,R0_data_188_4,R0_data_188_3,R0_data_188_2,
    R0_data_188_1,R0_data_188_0};
  wire [7:0] R0_data_189_0 = mem_189_0_R0_data;
  wire [7:0] R0_data_189_1 = mem_189_1_R0_data;
  wire [7:0] R0_data_189_2 = mem_189_2_R0_data;
  wire [7:0] R0_data_189_3 = mem_189_3_R0_data;
  wire [7:0] R0_data_189_4 = mem_189_4_R0_data;
  wire [7:0] R0_data_189_5 = mem_189_5_R0_data;
  wire [7:0] R0_data_189_6 = mem_189_6_R0_data;
  wire [7:0] R0_data_189_7 = mem_189_7_R0_data;
  wire [63:0] R0_data_189 = {R0_data_189_7,R0_data_189_6,R0_data_189_5,R0_data_189_4,R0_data_189_3,R0_data_189_2,
    R0_data_189_1,R0_data_189_0};
  wire [7:0] R0_data_190_0 = mem_190_0_R0_data;
  wire [7:0] R0_data_190_1 = mem_190_1_R0_data;
  wire [7:0] R0_data_190_2 = mem_190_2_R0_data;
  wire [7:0] R0_data_190_3 = mem_190_3_R0_data;
  wire [7:0] R0_data_190_4 = mem_190_4_R0_data;
  wire [7:0] R0_data_190_5 = mem_190_5_R0_data;
  wire [7:0] R0_data_190_6 = mem_190_6_R0_data;
  wire [7:0] R0_data_190_7 = mem_190_7_R0_data;
  wire [63:0] R0_data_190 = {R0_data_190_7,R0_data_190_6,R0_data_190_5,R0_data_190_4,R0_data_190_3,R0_data_190_2,
    R0_data_190_1,R0_data_190_0};
  wire [7:0] R0_data_191_0 = mem_191_0_R0_data;
  wire [7:0] R0_data_191_1 = mem_191_1_R0_data;
  wire [7:0] R0_data_191_2 = mem_191_2_R0_data;
  wire [7:0] R0_data_191_3 = mem_191_3_R0_data;
  wire [7:0] R0_data_191_4 = mem_191_4_R0_data;
  wire [7:0] R0_data_191_5 = mem_191_5_R0_data;
  wire [7:0] R0_data_191_6 = mem_191_6_R0_data;
  wire [7:0] R0_data_191_7 = mem_191_7_R0_data;
  wire [63:0] R0_data_191 = {R0_data_191_7,R0_data_191_6,R0_data_191_5,R0_data_191_4,R0_data_191_3,R0_data_191_2,
    R0_data_191_1,R0_data_191_0};
  wire [7:0] R0_data_192_0 = mem_192_0_R0_data;
  wire [7:0] R0_data_192_1 = mem_192_1_R0_data;
  wire [7:0] R0_data_192_2 = mem_192_2_R0_data;
  wire [7:0] R0_data_192_3 = mem_192_3_R0_data;
  wire [7:0] R0_data_192_4 = mem_192_4_R0_data;
  wire [7:0] R0_data_192_5 = mem_192_5_R0_data;
  wire [7:0] R0_data_192_6 = mem_192_6_R0_data;
  wire [7:0] R0_data_192_7 = mem_192_7_R0_data;
  wire [63:0] R0_data_192 = {R0_data_192_7,R0_data_192_6,R0_data_192_5,R0_data_192_4,R0_data_192_3,R0_data_192_2,
    R0_data_192_1,R0_data_192_0};
  wire [7:0] R0_data_193_0 = mem_193_0_R0_data;
  wire [7:0] R0_data_193_1 = mem_193_1_R0_data;
  wire [7:0] R0_data_193_2 = mem_193_2_R0_data;
  wire [7:0] R0_data_193_3 = mem_193_3_R0_data;
  wire [7:0] R0_data_193_4 = mem_193_4_R0_data;
  wire [7:0] R0_data_193_5 = mem_193_5_R0_data;
  wire [7:0] R0_data_193_6 = mem_193_6_R0_data;
  wire [7:0] R0_data_193_7 = mem_193_7_R0_data;
  wire [63:0] R0_data_193 = {R0_data_193_7,R0_data_193_6,R0_data_193_5,R0_data_193_4,R0_data_193_3,R0_data_193_2,
    R0_data_193_1,R0_data_193_0};
  wire [7:0] R0_data_194_0 = mem_194_0_R0_data;
  wire [7:0] R0_data_194_1 = mem_194_1_R0_data;
  wire [7:0] R0_data_194_2 = mem_194_2_R0_data;
  wire [7:0] R0_data_194_3 = mem_194_3_R0_data;
  wire [7:0] R0_data_194_4 = mem_194_4_R0_data;
  wire [7:0] R0_data_194_5 = mem_194_5_R0_data;
  wire [7:0] R0_data_194_6 = mem_194_6_R0_data;
  wire [7:0] R0_data_194_7 = mem_194_7_R0_data;
  wire [63:0] R0_data_194 = {R0_data_194_7,R0_data_194_6,R0_data_194_5,R0_data_194_4,R0_data_194_3,R0_data_194_2,
    R0_data_194_1,R0_data_194_0};
  wire [7:0] R0_data_195_0 = mem_195_0_R0_data;
  wire [7:0] R0_data_195_1 = mem_195_1_R0_data;
  wire [7:0] R0_data_195_2 = mem_195_2_R0_data;
  wire [7:0] R0_data_195_3 = mem_195_3_R0_data;
  wire [7:0] R0_data_195_4 = mem_195_4_R0_data;
  wire [7:0] R0_data_195_5 = mem_195_5_R0_data;
  wire [7:0] R0_data_195_6 = mem_195_6_R0_data;
  wire [7:0] R0_data_195_7 = mem_195_7_R0_data;
  wire [63:0] R0_data_195 = {R0_data_195_7,R0_data_195_6,R0_data_195_5,R0_data_195_4,R0_data_195_3,R0_data_195_2,
    R0_data_195_1,R0_data_195_0};
  wire [7:0] R0_data_196_0 = mem_196_0_R0_data;
  wire [7:0] R0_data_196_1 = mem_196_1_R0_data;
  wire [7:0] R0_data_196_2 = mem_196_2_R0_data;
  wire [7:0] R0_data_196_3 = mem_196_3_R0_data;
  wire [7:0] R0_data_196_4 = mem_196_4_R0_data;
  wire [7:0] R0_data_196_5 = mem_196_5_R0_data;
  wire [7:0] R0_data_196_6 = mem_196_6_R0_data;
  wire [7:0] R0_data_196_7 = mem_196_7_R0_data;
  wire [63:0] R0_data_196 = {R0_data_196_7,R0_data_196_6,R0_data_196_5,R0_data_196_4,R0_data_196_3,R0_data_196_2,
    R0_data_196_1,R0_data_196_0};
  wire [7:0] R0_data_197_0 = mem_197_0_R0_data;
  wire [7:0] R0_data_197_1 = mem_197_1_R0_data;
  wire [7:0] R0_data_197_2 = mem_197_2_R0_data;
  wire [7:0] R0_data_197_3 = mem_197_3_R0_data;
  wire [7:0] R0_data_197_4 = mem_197_4_R0_data;
  wire [7:0] R0_data_197_5 = mem_197_5_R0_data;
  wire [7:0] R0_data_197_6 = mem_197_6_R0_data;
  wire [7:0] R0_data_197_7 = mem_197_7_R0_data;
  wire [63:0] R0_data_197 = {R0_data_197_7,R0_data_197_6,R0_data_197_5,R0_data_197_4,R0_data_197_3,R0_data_197_2,
    R0_data_197_1,R0_data_197_0};
  wire [7:0] R0_data_198_0 = mem_198_0_R0_data;
  wire [7:0] R0_data_198_1 = mem_198_1_R0_data;
  wire [7:0] R0_data_198_2 = mem_198_2_R0_data;
  wire [7:0] R0_data_198_3 = mem_198_3_R0_data;
  wire [7:0] R0_data_198_4 = mem_198_4_R0_data;
  wire [7:0] R0_data_198_5 = mem_198_5_R0_data;
  wire [7:0] R0_data_198_6 = mem_198_6_R0_data;
  wire [7:0] R0_data_198_7 = mem_198_7_R0_data;
  wire [63:0] R0_data_198 = {R0_data_198_7,R0_data_198_6,R0_data_198_5,R0_data_198_4,R0_data_198_3,R0_data_198_2,
    R0_data_198_1,R0_data_198_0};
  wire [7:0] R0_data_199_0 = mem_199_0_R0_data;
  wire [7:0] R0_data_199_1 = mem_199_1_R0_data;
  wire [7:0] R0_data_199_2 = mem_199_2_R0_data;
  wire [7:0] R0_data_199_3 = mem_199_3_R0_data;
  wire [7:0] R0_data_199_4 = mem_199_4_R0_data;
  wire [7:0] R0_data_199_5 = mem_199_5_R0_data;
  wire [7:0] R0_data_199_6 = mem_199_6_R0_data;
  wire [7:0] R0_data_199_7 = mem_199_7_R0_data;
  wire [63:0] R0_data_199 = {R0_data_199_7,R0_data_199_6,R0_data_199_5,R0_data_199_4,R0_data_199_3,R0_data_199_2,
    R0_data_199_1,R0_data_199_0};
  wire [7:0] R0_data_200_0 = mem_200_0_R0_data;
  wire [7:0] R0_data_200_1 = mem_200_1_R0_data;
  wire [7:0] R0_data_200_2 = mem_200_2_R0_data;
  wire [7:0] R0_data_200_3 = mem_200_3_R0_data;
  wire [7:0] R0_data_200_4 = mem_200_4_R0_data;
  wire [7:0] R0_data_200_5 = mem_200_5_R0_data;
  wire [7:0] R0_data_200_6 = mem_200_6_R0_data;
  wire [7:0] R0_data_200_7 = mem_200_7_R0_data;
  wire [63:0] R0_data_200 = {R0_data_200_7,R0_data_200_6,R0_data_200_5,R0_data_200_4,R0_data_200_3,R0_data_200_2,
    R0_data_200_1,R0_data_200_0};
  wire [7:0] R0_data_201_0 = mem_201_0_R0_data;
  wire [7:0] R0_data_201_1 = mem_201_1_R0_data;
  wire [7:0] R0_data_201_2 = mem_201_2_R0_data;
  wire [7:0] R0_data_201_3 = mem_201_3_R0_data;
  wire [7:0] R0_data_201_4 = mem_201_4_R0_data;
  wire [7:0] R0_data_201_5 = mem_201_5_R0_data;
  wire [7:0] R0_data_201_6 = mem_201_6_R0_data;
  wire [7:0] R0_data_201_7 = mem_201_7_R0_data;
  wire [63:0] R0_data_201 = {R0_data_201_7,R0_data_201_6,R0_data_201_5,R0_data_201_4,R0_data_201_3,R0_data_201_2,
    R0_data_201_1,R0_data_201_0};
  wire [7:0] R0_data_202_0 = mem_202_0_R0_data;
  wire [7:0] R0_data_202_1 = mem_202_1_R0_data;
  wire [7:0] R0_data_202_2 = mem_202_2_R0_data;
  wire [7:0] R0_data_202_3 = mem_202_3_R0_data;
  wire [7:0] R0_data_202_4 = mem_202_4_R0_data;
  wire [7:0] R0_data_202_5 = mem_202_5_R0_data;
  wire [7:0] R0_data_202_6 = mem_202_6_R0_data;
  wire [7:0] R0_data_202_7 = mem_202_7_R0_data;
  wire [63:0] R0_data_202 = {R0_data_202_7,R0_data_202_6,R0_data_202_5,R0_data_202_4,R0_data_202_3,R0_data_202_2,
    R0_data_202_1,R0_data_202_0};
  wire [7:0] R0_data_203_0 = mem_203_0_R0_data;
  wire [7:0] R0_data_203_1 = mem_203_1_R0_data;
  wire [7:0] R0_data_203_2 = mem_203_2_R0_data;
  wire [7:0] R0_data_203_3 = mem_203_3_R0_data;
  wire [7:0] R0_data_203_4 = mem_203_4_R0_data;
  wire [7:0] R0_data_203_5 = mem_203_5_R0_data;
  wire [7:0] R0_data_203_6 = mem_203_6_R0_data;
  wire [7:0] R0_data_203_7 = mem_203_7_R0_data;
  wire [63:0] R0_data_203 = {R0_data_203_7,R0_data_203_6,R0_data_203_5,R0_data_203_4,R0_data_203_3,R0_data_203_2,
    R0_data_203_1,R0_data_203_0};
  wire [7:0] R0_data_204_0 = mem_204_0_R0_data;
  wire [7:0] R0_data_204_1 = mem_204_1_R0_data;
  wire [7:0] R0_data_204_2 = mem_204_2_R0_data;
  wire [7:0] R0_data_204_3 = mem_204_3_R0_data;
  wire [7:0] R0_data_204_4 = mem_204_4_R0_data;
  wire [7:0] R0_data_204_5 = mem_204_5_R0_data;
  wire [7:0] R0_data_204_6 = mem_204_6_R0_data;
  wire [7:0] R0_data_204_7 = mem_204_7_R0_data;
  wire [63:0] R0_data_204 = {R0_data_204_7,R0_data_204_6,R0_data_204_5,R0_data_204_4,R0_data_204_3,R0_data_204_2,
    R0_data_204_1,R0_data_204_0};
  wire [7:0] R0_data_205_0 = mem_205_0_R0_data;
  wire [7:0] R0_data_205_1 = mem_205_1_R0_data;
  wire [7:0] R0_data_205_2 = mem_205_2_R0_data;
  wire [7:0] R0_data_205_3 = mem_205_3_R0_data;
  wire [7:0] R0_data_205_4 = mem_205_4_R0_data;
  wire [7:0] R0_data_205_5 = mem_205_5_R0_data;
  wire [7:0] R0_data_205_6 = mem_205_6_R0_data;
  wire [7:0] R0_data_205_7 = mem_205_7_R0_data;
  wire [63:0] R0_data_205 = {R0_data_205_7,R0_data_205_6,R0_data_205_5,R0_data_205_4,R0_data_205_3,R0_data_205_2,
    R0_data_205_1,R0_data_205_0};
  wire [7:0] R0_data_206_0 = mem_206_0_R0_data;
  wire [7:0] R0_data_206_1 = mem_206_1_R0_data;
  wire [7:0] R0_data_206_2 = mem_206_2_R0_data;
  wire [7:0] R0_data_206_3 = mem_206_3_R0_data;
  wire [7:0] R0_data_206_4 = mem_206_4_R0_data;
  wire [7:0] R0_data_206_5 = mem_206_5_R0_data;
  wire [7:0] R0_data_206_6 = mem_206_6_R0_data;
  wire [7:0] R0_data_206_7 = mem_206_7_R0_data;
  wire [63:0] R0_data_206 = {R0_data_206_7,R0_data_206_6,R0_data_206_5,R0_data_206_4,R0_data_206_3,R0_data_206_2,
    R0_data_206_1,R0_data_206_0};
  wire [7:0] R0_data_207_0 = mem_207_0_R0_data;
  wire [7:0] R0_data_207_1 = mem_207_1_R0_data;
  wire [7:0] R0_data_207_2 = mem_207_2_R0_data;
  wire [7:0] R0_data_207_3 = mem_207_3_R0_data;
  wire [7:0] R0_data_207_4 = mem_207_4_R0_data;
  wire [7:0] R0_data_207_5 = mem_207_5_R0_data;
  wire [7:0] R0_data_207_6 = mem_207_6_R0_data;
  wire [7:0] R0_data_207_7 = mem_207_7_R0_data;
  wire [63:0] R0_data_207 = {R0_data_207_7,R0_data_207_6,R0_data_207_5,R0_data_207_4,R0_data_207_3,R0_data_207_2,
    R0_data_207_1,R0_data_207_0};
  wire [7:0] R0_data_208_0 = mem_208_0_R0_data;
  wire [7:0] R0_data_208_1 = mem_208_1_R0_data;
  wire [7:0] R0_data_208_2 = mem_208_2_R0_data;
  wire [7:0] R0_data_208_3 = mem_208_3_R0_data;
  wire [7:0] R0_data_208_4 = mem_208_4_R0_data;
  wire [7:0] R0_data_208_5 = mem_208_5_R0_data;
  wire [7:0] R0_data_208_6 = mem_208_6_R0_data;
  wire [7:0] R0_data_208_7 = mem_208_7_R0_data;
  wire [63:0] R0_data_208 = {R0_data_208_7,R0_data_208_6,R0_data_208_5,R0_data_208_4,R0_data_208_3,R0_data_208_2,
    R0_data_208_1,R0_data_208_0};
  wire [7:0] R0_data_209_0 = mem_209_0_R0_data;
  wire [7:0] R0_data_209_1 = mem_209_1_R0_data;
  wire [7:0] R0_data_209_2 = mem_209_2_R0_data;
  wire [7:0] R0_data_209_3 = mem_209_3_R0_data;
  wire [7:0] R0_data_209_4 = mem_209_4_R0_data;
  wire [7:0] R0_data_209_5 = mem_209_5_R0_data;
  wire [7:0] R0_data_209_6 = mem_209_6_R0_data;
  wire [7:0] R0_data_209_7 = mem_209_7_R0_data;
  wire [63:0] R0_data_209 = {R0_data_209_7,R0_data_209_6,R0_data_209_5,R0_data_209_4,R0_data_209_3,R0_data_209_2,
    R0_data_209_1,R0_data_209_0};
  wire [7:0] R0_data_210_0 = mem_210_0_R0_data;
  wire [7:0] R0_data_210_1 = mem_210_1_R0_data;
  wire [7:0] R0_data_210_2 = mem_210_2_R0_data;
  wire [7:0] R0_data_210_3 = mem_210_3_R0_data;
  wire [7:0] R0_data_210_4 = mem_210_4_R0_data;
  wire [7:0] R0_data_210_5 = mem_210_5_R0_data;
  wire [7:0] R0_data_210_6 = mem_210_6_R0_data;
  wire [7:0] R0_data_210_7 = mem_210_7_R0_data;
  wire [63:0] R0_data_210 = {R0_data_210_7,R0_data_210_6,R0_data_210_5,R0_data_210_4,R0_data_210_3,R0_data_210_2,
    R0_data_210_1,R0_data_210_0};
  wire [7:0] R0_data_211_0 = mem_211_0_R0_data;
  wire [7:0] R0_data_211_1 = mem_211_1_R0_data;
  wire [7:0] R0_data_211_2 = mem_211_2_R0_data;
  wire [7:0] R0_data_211_3 = mem_211_3_R0_data;
  wire [7:0] R0_data_211_4 = mem_211_4_R0_data;
  wire [7:0] R0_data_211_5 = mem_211_5_R0_data;
  wire [7:0] R0_data_211_6 = mem_211_6_R0_data;
  wire [7:0] R0_data_211_7 = mem_211_7_R0_data;
  wire [63:0] R0_data_211 = {R0_data_211_7,R0_data_211_6,R0_data_211_5,R0_data_211_4,R0_data_211_3,R0_data_211_2,
    R0_data_211_1,R0_data_211_0};
  wire [7:0] R0_data_212_0 = mem_212_0_R0_data;
  wire [7:0] R0_data_212_1 = mem_212_1_R0_data;
  wire [7:0] R0_data_212_2 = mem_212_2_R0_data;
  wire [7:0] R0_data_212_3 = mem_212_3_R0_data;
  wire [7:0] R0_data_212_4 = mem_212_4_R0_data;
  wire [7:0] R0_data_212_5 = mem_212_5_R0_data;
  wire [7:0] R0_data_212_6 = mem_212_6_R0_data;
  wire [7:0] R0_data_212_7 = mem_212_7_R0_data;
  wire [63:0] R0_data_212 = {R0_data_212_7,R0_data_212_6,R0_data_212_5,R0_data_212_4,R0_data_212_3,R0_data_212_2,
    R0_data_212_1,R0_data_212_0};
  wire [7:0] R0_data_213_0 = mem_213_0_R0_data;
  wire [7:0] R0_data_213_1 = mem_213_1_R0_data;
  wire [7:0] R0_data_213_2 = mem_213_2_R0_data;
  wire [7:0] R0_data_213_3 = mem_213_3_R0_data;
  wire [7:0] R0_data_213_4 = mem_213_4_R0_data;
  wire [7:0] R0_data_213_5 = mem_213_5_R0_data;
  wire [7:0] R0_data_213_6 = mem_213_6_R0_data;
  wire [7:0] R0_data_213_7 = mem_213_7_R0_data;
  wire [63:0] R0_data_213 = {R0_data_213_7,R0_data_213_6,R0_data_213_5,R0_data_213_4,R0_data_213_3,R0_data_213_2,
    R0_data_213_1,R0_data_213_0};
  wire [7:0] R0_data_214_0 = mem_214_0_R0_data;
  wire [7:0] R0_data_214_1 = mem_214_1_R0_data;
  wire [7:0] R0_data_214_2 = mem_214_2_R0_data;
  wire [7:0] R0_data_214_3 = mem_214_3_R0_data;
  wire [7:0] R0_data_214_4 = mem_214_4_R0_data;
  wire [7:0] R0_data_214_5 = mem_214_5_R0_data;
  wire [7:0] R0_data_214_6 = mem_214_6_R0_data;
  wire [7:0] R0_data_214_7 = mem_214_7_R0_data;
  wire [63:0] R0_data_214 = {R0_data_214_7,R0_data_214_6,R0_data_214_5,R0_data_214_4,R0_data_214_3,R0_data_214_2,
    R0_data_214_1,R0_data_214_0};
  wire [7:0] R0_data_215_0 = mem_215_0_R0_data;
  wire [7:0] R0_data_215_1 = mem_215_1_R0_data;
  wire [7:0] R0_data_215_2 = mem_215_2_R0_data;
  wire [7:0] R0_data_215_3 = mem_215_3_R0_data;
  wire [7:0] R0_data_215_4 = mem_215_4_R0_data;
  wire [7:0] R0_data_215_5 = mem_215_5_R0_data;
  wire [7:0] R0_data_215_6 = mem_215_6_R0_data;
  wire [7:0] R0_data_215_7 = mem_215_7_R0_data;
  wire [63:0] R0_data_215 = {R0_data_215_7,R0_data_215_6,R0_data_215_5,R0_data_215_4,R0_data_215_3,R0_data_215_2,
    R0_data_215_1,R0_data_215_0};
  wire [7:0] R0_data_216_0 = mem_216_0_R0_data;
  wire [7:0] R0_data_216_1 = mem_216_1_R0_data;
  wire [7:0] R0_data_216_2 = mem_216_2_R0_data;
  wire [7:0] R0_data_216_3 = mem_216_3_R0_data;
  wire [7:0] R0_data_216_4 = mem_216_4_R0_data;
  wire [7:0] R0_data_216_5 = mem_216_5_R0_data;
  wire [7:0] R0_data_216_6 = mem_216_6_R0_data;
  wire [7:0] R0_data_216_7 = mem_216_7_R0_data;
  wire [63:0] R0_data_216 = {R0_data_216_7,R0_data_216_6,R0_data_216_5,R0_data_216_4,R0_data_216_3,R0_data_216_2,
    R0_data_216_1,R0_data_216_0};
  wire [7:0] R0_data_217_0 = mem_217_0_R0_data;
  wire [7:0] R0_data_217_1 = mem_217_1_R0_data;
  wire [7:0] R0_data_217_2 = mem_217_2_R0_data;
  wire [7:0] R0_data_217_3 = mem_217_3_R0_data;
  wire [7:0] R0_data_217_4 = mem_217_4_R0_data;
  wire [7:0] R0_data_217_5 = mem_217_5_R0_data;
  wire [7:0] R0_data_217_6 = mem_217_6_R0_data;
  wire [7:0] R0_data_217_7 = mem_217_7_R0_data;
  wire [63:0] R0_data_217 = {R0_data_217_7,R0_data_217_6,R0_data_217_5,R0_data_217_4,R0_data_217_3,R0_data_217_2,
    R0_data_217_1,R0_data_217_0};
  wire [7:0] R0_data_218_0 = mem_218_0_R0_data;
  wire [7:0] R0_data_218_1 = mem_218_1_R0_data;
  wire [7:0] R0_data_218_2 = mem_218_2_R0_data;
  wire [7:0] R0_data_218_3 = mem_218_3_R0_data;
  wire [7:0] R0_data_218_4 = mem_218_4_R0_data;
  wire [7:0] R0_data_218_5 = mem_218_5_R0_data;
  wire [7:0] R0_data_218_6 = mem_218_6_R0_data;
  wire [7:0] R0_data_218_7 = mem_218_7_R0_data;
  wire [63:0] R0_data_218 = {R0_data_218_7,R0_data_218_6,R0_data_218_5,R0_data_218_4,R0_data_218_3,R0_data_218_2,
    R0_data_218_1,R0_data_218_0};
  wire [7:0] R0_data_219_0 = mem_219_0_R0_data;
  wire [7:0] R0_data_219_1 = mem_219_1_R0_data;
  wire [7:0] R0_data_219_2 = mem_219_2_R0_data;
  wire [7:0] R0_data_219_3 = mem_219_3_R0_data;
  wire [7:0] R0_data_219_4 = mem_219_4_R0_data;
  wire [7:0] R0_data_219_5 = mem_219_5_R0_data;
  wire [7:0] R0_data_219_6 = mem_219_6_R0_data;
  wire [7:0] R0_data_219_7 = mem_219_7_R0_data;
  wire [63:0] R0_data_219 = {R0_data_219_7,R0_data_219_6,R0_data_219_5,R0_data_219_4,R0_data_219_3,R0_data_219_2,
    R0_data_219_1,R0_data_219_0};
  wire [7:0] R0_data_220_0 = mem_220_0_R0_data;
  wire [7:0] R0_data_220_1 = mem_220_1_R0_data;
  wire [7:0] R0_data_220_2 = mem_220_2_R0_data;
  wire [7:0] R0_data_220_3 = mem_220_3_R0_data;
  wire [7:0] R0_data_220_4 = mem_220_4_R0_data;
  wire [7:0] R0_data_220_5 = mem_220_5_R0_data;
  wire [7:0] R0_data_220_6 = mem_220_6_R0_data;
  wire [7:0] R0_data_220_7 = mem_220_7_R0_data;
  wire [63:0] R0_data_220 = {R0_data_220_7,R0_data_220_6,R0_data_220_5,R0_data_220_4,R0_data_220_3,R0_data_220_2,
    R0_data_220_1,R0_data_220_0};
  wire [7:0] R0_data_221_0 = mem_221_0_R0_data;
  wire [7:0] R0_data_221_1 = mem_221_1_R0_data;
  wire [7:0] R0_data_221_2 = mem_221_2_R0_data;
  wire [7:0] R0_data_221_3 = mem_221_3_R0_data;
  wire [7:0] R0_data_221_4 = mem_221_4_R0_data;
  wire [7:0] R0_data_221_5 = mem_221_5_R0_data;
  wire [7:0] R0_data_221_6 = mem_221_6_R0_data;
  wire [7:0] R0_data_221_7 = mem_221_7_R0_data;
  wire [63:0] R0_data_221 = {R0_data_221_7,R0_data_221_6,R0_data_221_5,R0_data_221_4,R0_data_221_3,R0_data_221_2,
    R0_data_221_1,R0_data_221_0};
  wire [7:0] R0_data_222_0 = mem_222_0_R0_data;
  wire [7:0] R0_data_222_1 = mem_222_1_R0_data;
  wire [7:0] R0_data_222_2 = mem_222_2_R0_data;
  wire [7:0] R0_data_222_3 = mem_222_3_R0_data;
  wire [7:0] R0_data_222_4 = mem_222_4_R0_data;
  wire [7:0] R0_data_222_5 = mem_222_5_R0_data;
  wire [7:0] R0_data_222_6 = mem_222_6_R0_data;
  wire [7:0] R0_data_222_7 = mem_222_7_R0_data;
  wire [63:0] R0_data_222 = {R0_data_222_7,R0_data_222_6,R0_data_222_5,R0_data_222_4,R0_data_222_3,R0_data_222_2,
    R0_data_222_1,R0_data_222_0};
  wire [7:0] R0_data_223_0 = mem_223_0_R0_data;
  wire [7:0] R0_data_223_1 = mem_223_1_R0_data;
  wire [7:0] R0_data_223_2 = mem_223_2_R0_data;
  wire [7:0] R0_data_223_3 = mem_223_3_R0_data;
  wire [7:0] R0_data_223_4 = mem_223_4_R0_data;
  wire [7:0] R0_data_223_5 = mem_223_5_R0_data;
  wire [7:0] R0_data_223_6 = mem_223_6_R0_data;
  wire [7:0] R0_data_223_7 = mem_223_7_R0_data;
  wire [63:0] R0_data_223 = {R0_data_223_7,R0_data_223_6,R0_data_223_5,R0_data_223_4,R0_data_223_3,R0_data_223_2,
    R0_data_223_1,R0_data_223_0};
  wire [7:0] R0_data_224_0 = mem_224_0_R0_data;
  wire [7:0] R0_data_224_1 = mem_224_1_R0_data;
  wire [7:0] R0_data_224_2 = mem_224_2_R0_data;
  wire [7:0] R0_data_224_3 = mem_224_3_R0_data;
  wire [7:0] R0_data_224_4 = mem_224_4_R0_data;
  wire [7:0] R0_data_224_5 = mem_224_5_R0_data;
  wire [7:0] R0_data_224_6 = mem_224_6_R0_data;
  wire [7:0] R0_data_224_7 = mem_224_7_R0_data;
  wire [63:0] R0_data_224 = {R0_data_224_7,R0_data_224_6,R0_data_224_5,R0_data_224_4,R0_data_224_3,R0_data_224_2,
    R0_data_224_1,R0_data_224_0};
  wire [7:0] R0_data_225_0 = mem_225_0_R0_data;
  wire [7:0] R0_data_225_1 = mem_225_1_R0_data;
  wire [7:0] R0_data_225_2 = mem_225_2_R0_data;
  wire [7:0] R0_data_225_3 = mem_225_3_R0_data;
  wire [7:0] R0_data_225_4 = mem_225_4_R0_data;
  wire [7:0] R0_data_225_5 = mem_225_5_R0_data;
  wire [7:0] R0_data_225_6 = mem_225_6_R0_data;
  wire [7:0] R0_data_225_7 = mem_225_7_R0_data;
  wire [63:0] R0_data_225 = {R0_data_225_7,R0_data_225_6,R0_data_225_5,R0_data_225_4,R0_data_225_3,R0_data_225_2,
    R0_data_225_1,R0_data_225_0};
  wire [7:0] R0_data_226_0 = mem_226_0_R0_data;
  wire [7:0] R0_data_226_1 = mem_226_1_R0_data;
  wire [7:0] R0_data_226_2 = mem_226_2_R0_data;
  wire [7:0] R0_data_226_3 = mem_226_3_R0_data;
  wire [7:0] R0_data_226_4 = mem_226_4_R0_data;
  wire [7:0] R0_data_226_5 = mem_226_5_R0_data;
  wire [7:0] R0_data_226_6 = mem_226_6_R0_data;
  wire [7:0] R0_data_226_7 = mem_226_7_R0_data;
  wire [63:0] R0_data_226 = {R0_data_226_7,R0_data_226_6,R0_data_226_5,R0_data_226_4,R0_data_226_3,R0_data_226_2,
    R0_data_226_1,R0_data_226_0};
  wire [7:0] R0_data_227_0 = mem_227_0_R0_data;
  wire [7:0] R0_data_227_1 = mem_227_1_R0_data;
  wire [7:0] R0_data_227_2 = mem_227_2_R0_data;
  wire [7:0] R0_data_227_3 = mem_227_3_R0_data;
  wire [7:0] R0_data_227_4 = mem_227_4_R0_data;
  wire [7:0] R0_data_227_5 = mem_227_5_R0_data;
  wire [7:0] R0_data_227_6 = mem_227_6_R0_data;
  wire [7:0] R0_data_227_7 = mem_227_7_R0_data;
  wire [63:0] R0_data_227 = {R0_data_227_7,R0_data_227_6,R0_data_227_5,R0_data_227_4,R0_data_227_3,R0_data_227_2,
    R0_data_227_1,R0_data_227_0};
  wire [7:0] R0_data_228_0 = mem_228_0_R0_data;
  wire [7:0] R0_data_228_1 = mem_228_1_R0_data;
  wire [7:0] R0_data_228_2 = mem_228_2_R0_data;
  wire [7:0] R0_data_228_3 = mem_228_3_R0_data;
  wire [7:0] R0_data_228_4 = mem_228_4_R0_data;
  wire [7:0] R0_data_228_5 = mem_228_5_R0_data;
  wire [7:0] R0_data_228_6 = mem_228_6_R0_data;
  wire [7:0] R0_data_228_7 = mem_228_7_R0_data;
  wire [63:0] R0_data_228 = {R0_data_228_7,R0_data_228_6,R0_data_228_5,R0_data_228_4,R0_data_228_3,R0_data_228_2,
    R0_data_228_1,R0_data_228_0};
  wire [7:0] R0_data_229_0 = mem_229_0_R0_data;
  wire [7:0] R0_data_229_1 = mem_229_1_R0_data;
  wire [7:0] R0_data_229_2 = mem_229_2_R0_data;
  wire [7:0] R0_data_229_3 = mem_229_3_R0_data;
  wire [7:0] R0_data_229_4 = mem_229_4_R0_data;
  wire [7:0] R0_data_229_5 = mem_229_5_R0_data;
  wire [7:0] R0_data_229_6 = mem_229_6_R0_data;
  wire [7:0] R0_data_229_7 = mem_229_7_R0_data;
  wire [63:0] R0_data_229 = {R0_data_229_7,R0_data_229_6,R0_data_229_5,R0_data_229_4,R0_data_229_3,R0_data_229_2,
    R0_data_229_1,R0_data_229_0};
  wire [7:0] R0_data_230_0 = mem_230_0_R0_data;
  wire [7:0] R0_data_230_1 = mem_230_1_R0_data;
  wire [7:0] R0_data_230_2 = mem_230_2_R0_data;
  wire [7:0] R0_data_230_3 = mem_230_3_R0_data;
  wire [7:0] R0_data_230_4 = mem_230_4_R0_data;
  wire [7:0] R0_data_230_5 = mem_230_5_R0_data;
  wire [7:0] R0_data_230_6 = mem_230_6_R0_data;
  wire [7:0] R0_data_230_7 = mem_230_7_R0_data;
  wire [63:0] R0_data_230 = {R0_data_230_7,R0_data_230_6,R0_data_230_5,R0_data_230_4,R0_data_230_3,R0_data_230_2,
    R0_data_230_1,R0_data_230_0};
  wire [7:0] R0_data_231_0 = mem_231_0_R0_data;
  wire [7:0] R0_data_231_1 = mem_231_1_R0_data;
  wire [7:0] R0_data_231_2 = mem_231_2_R0_data;
  wire [7:0] R0_data_231_3 = mem_231_3_R0_data;
  wire [7:0] R0_data_231_4 = mem_231_4_R0_data;
  wire [7:0] R0_data_231_5 = mem_231_5_R0_data;
  wire [7:0] R0_data_231_6 = mem_231_6_R0_data;
  wire [7:0] R0_data_231_7 = mem_231_7_R0_data;
  wire [63:0] R0_data_231 = {R0_data_231_7,R0_data_231_6,R0_data_231_5,R0_data_231_4,R0_data_231_3,R0_data_231_2,
    R0_data_231_1,R0_data_231_0};
  wire [7:0] R0_data_232_0 = mem_232_0_R0_data;
  wire [7:0] R0_data_232_1 = mem_232_1_R0_data;
  wire [7:0] R0_data_232_2 = mem_232_2_R0_data;
  wire [7:0] R0_data_232_3 = mem_232_3_R0_data;
  wire [7:0] R0_data_232_4 = mem_232_4_R0_data;
  wire [7:0] R0_data_232_5 = mem_232_5_R0_data;
  wire [7:0] R0_data_232_6 = mem_232_6_R0_data;
  wire [7:0] R0_data_232_7 = mem_232_7_R0_data;
  wire [63:0] R0_data_232 = {R0_data_232_7,R0_data_232_6,R0_data_232_5,R0_data_232_4,R0_data_232_3,R0_data_232_2,
    R0_data_232_1,R0_data_232_0};
  wire [7:0] R0_data_233_0 = mem_233_0_R0_data;
  wire [7:0] R0_data_233_1 = mem_233_1_R0_data;
  wire [7:0] R0_data_233_2 = mem_233_2_R0_data;
  wire [7:0] R0_data_233_3 = mem_233_3_R0_data;
  wire [7:0] R0_data_233_4 = mem_233_4_R0_data;
  wire [7:0] R0_data_233_5 = mem_233_5_R0_data;
  wire [7:0] R0_data_233_6 = mem_233_6_R0_data;
  wire [7:0] R0_data_233_7 = mem_233_7_R0_data;
  wire [63:0] R0_data_233 = {R0_data_233_7,R0_data_233_6,R0_data_233_5,R0_data_233_4,R0_data_233_3,R0_data_233_2,
    R0_data_233_1,R0_data_233_0};
  wire [7:0] R0_data_234_0 = mem_234_0_R0_data;
  wire [7:0] R0_data_234_1 = mem_234_1_R0_data;
  wire [7:0] R0_data_234_2 = mem_234_2_R0_data;
  wire [7:0] R0_data_234_3 = mem_234_3_R0_data;
  wire [7:0] R0_data_234_4 = mem_234_4_R0_data;
  wire [7:0] R0_data_234_5 = mem_234_5_R0_data;
  wire [7:0] R0_data_234_6 = mem_234_6_R0_data;
  wire [7:0] R0_data_234_7 = mem_234_7_R0_data;
  wire [63:0] R0_data_234 = {R0_data_234_7,R0_data_234_6,R0_data_234_5,R0_data_234_4,R0_data_234_3,R0_data_234_2,
    R0_data_234_1,R0_data_234_0};
  wire [7:0] R0_data_235_0 = mem_235_0_R0_data;
  wire [7:0] R0_data_235_1 = mem_235_1_R0_data;
  wire [7:0] R0_data_235_2 = mem_235_2_R0_data;
  wire [7:0] R0_data_235_3 = mem_235_3_R0_data;
  wire [7:0] R0_data_235_4 = mem_235_4_R0_data;
  wire [7:0] R0_data_235_5 = mem_235_5_R0_data;
  wire [7:0] R0_data_235_6 = mem_235_6_R0_data;
  wire [7:0] R0_data_235_7 = mem_235_7_R0_data;
  wire [63:0] R0_data_235 = {R0_data_235_7,R0_data_235_6,R0_data_235_5,R0_data_235_4,R0_data_235_3,R0_data_235_2,
    R0_data_235_1,R0_data_235_0};
  wire [7:0] R0_data_236_0 = mem_236_0_R0_data;
  wire [7:0] R0_data_236_1 = mem_236_1_R0_data;
  wire [7:0] R0_data_236_2 = mem_236_2_R0_data;
  wire [7:0] R0_data_236_3 = mem_236_3_R0_data;
  wire [7:0] R0_data_236_4 = mem_236_4_R0_data;
  wire [7:0] R0_data_236_5 = mem_236_5_R0_data;
  wire [7:0] R0_data_236_6 = mem_236_6_R0_data;
  wire [7:0] R0_data_236_7 = mem_236_7_R0_data;
  wire [63:0] R0_data_236 = {R0_data_236_7,R0_data_236_6,R0_data_236_5,R0_data_236_4,R0_data_236_3,R0_data_236_2,
    R0_data_236_1,R0_data_236_0};
  wire [7:0] R0_data_237_0 = mem_237_0_R0_data;
  wire [7:0] R0_data_237_1 = mem_237_1_R0_data;
  wire [7:0] R0_data_237_2 = mem_237_2_R0_data;
  wire [7:0] R0_data_237_3 = mem_237_3_R0_data;
  wire [7:0] R0_data_237_4 = mem_237_4_R0_data;
  wire [7:0] R0_data_237_5 = mem_237_5_R0_data;
  wire [7:0] R0_data_237_6 = mem_237_6_R0_data;
  wire [7:0] R0_data_237_7 = mem_237_7_R0_data;
  wire [63:0] R0_data_237 = {R0_data_237_7,R0_data_237_6,R0_data_237_5,R0_data_237_4,R0_data_237_3,R0_data_237_2,
    R0_data_237_1,R0_data_237_0};
  wire [7:0] R0_data_238_0 = mem_238_0_R0_data;
  wire [7:0] R0_data_238_1 = mem_238_1_R0_data;
  wire [7:0] R0_data_238_2 = mem_238_2_R0_data;
  wire [7:0] R0_data_238_3 = mem_238_3_R0_data;
  wire [7:0] R0_data_238_4 = mem_238_4_R0_data;
  wire [7:0] R0_data_238_5 = mem_238_5_R0_data;
  wire [7:0] R0_data_238_6 = mem_238_6_R0_data;
  wire [7:0] R0_data_238_7 = mem_238_7_R0_data;
  wire [63:0] R0_data_238 = {R0_data_238_7,R0_data_238_6,R0_data_238_5,R0_data_238_4,R0_data_238_3,R0_data_238_2,
    R0_data_238_1,R0_data_238_0};
  wire [7:0] R0_data_239_0 = mem_239_0_R0_data;
  wire [7:0] R0_data_239_1 = mem_239_1_R0_data;
  wire [7:0] R0_data_239_2 = mem_239_2_R0_data;
  wire [7:0] R0_data_239_3 = mem_239_3_R0_data;
  wire [7:0] R0_data_239_4 = mem_239_4_R0_data;
  wire [7:0] R0_data_239_5 = mem_239_5_R0_data;
  wire [7:0] R0_data_239_6 = mem_239_6_R0_data;
  wire [7:0] R0_data_239_7 = mem_239_7_R0_data;
  wire [63:0] R0_data_239 = {R0_data_239_7,R0_data_239_6,R0_data_239_5,R0_data_239_4,R0_data_239_3,R0_data_239_2,
    R0_data_239_1,R0_data_239_0};
  wire [7:0] R0_data_240_0 = mem_240_0_R0_data;
  wire [7:0] R0_data_240_1 = mem_240_1_R0_data;
  wire [7:0] R0_data_240_2 = mem_240_2_R0_data;
  wire [7:0] R0_data_240_3 = mem_240_3_R0_data;
  wire [7:0] R0_data_240_4 = mem_240_4_R0_data;
  wire [7:0] R0_data_240_5 = mem_240_5_R0_data;
  wire [7:0] R0_data_240_6 = mem_240_6_R0_data;
  wire [7:0] R0_data_240_7 = mem_240_7_R0_data;
  wire [63:0] R0_data_240 = {R0_data_240_7,R0_data_240_6,R0_data_240_5,R0_data_240_4,R0_data_240_3,R0_data_240_2,
    R0_data_240_1,R0_data_240_0};
  wire [7:0] R0_data_241_0 = mem_241_0_R0_data;
  wire [7:0] R0_data_241_1 = mem_241_1_R0_data;
  wire [7:0] R0_data_241_2 = mem_241_2_R0_data;
  wire [7:0] R0_data_241_3 = mem_241_3_R0_data;
  wire [7:0] R0_data_241_4 = mem_241_4_R0_data;
  wire [7:0] R0_data_241_5 = mem_241_5_R0_data;
  wire [7:0] R0_data_241_6 = mem_241_6_R0_data;
  wire [7:0] R0_data_241_7 = mem_241_7_R0_data;
  wire [63:0] R0_data_241 = {R0_data_241_7,R0_data_241_6,R0_data_241_5,R0_data_241_4,R0_data_241_3,R0_data_241_2,
    R0_data_241_1,R0_data_241_0};
  wire [7:0] R0_data_242_0 = mem_242_0_R0_data;
  wire [7:0] R0_data_242_1 = mem_242_1_R0_data;
  wire [7:0] R0_data_242_2 = mem_242_2_R0_data;
  wire [7:0] R0_data_242_3 = mem_242_3_R0_data;
  wire [7:0] R0_data_242_4 = mem_242_4_R0_data;
  wire [7:0] R0_data_242_5 = mem_242_5_R0_data;
  wire [7:0] R0_data_242_6 = mem_242_6_R0_data;
  wire [7:0] R0_data_242_7 = mem_242_7_R0_data;
  wire [63:0] R0_data_242 = {R0_data_242_7,R0_data_242_6,R0_data_242_5,R0_data_242_4,R0_data_242_3,R0_data_242_2,
    R0_data_242_1,R0_data_242_0};
  wire [7:0] R0_data_243_0 = mem_243_0_R0_data;
  wire [7:0] R0_data_243_1 = mem_243_1_R0_data;
  wire [7:0] R0_data_243_2 = mem_243_2_R0_data;
  wire [7:0] R0_data_243_3 = mem_243_3_R0_data;
  wire [7:0] R0_data_243_4 = mem_243_4_R0_data;
  wire [7:0] R0_data_243_5 = mem_243_5_R0_data;
  wire [7:0] R0_data_243_6 = mem_243_6_R0_data;
  wire [7:0] R0_data_243_7 = mem_243_7_R0_data;
  wire [63:0] R0_data_243 = {R0_data_243_7,R0_data_243_6,R0_data_243_5,R0_data_243_4,R0_data_243_3,R0_data_243_2,
    R0_data_243_1,R0_data_243_0};
  wire [7:0] R0_data_244_0 = mem_244_0_R0_data;
  wire [7:0] R0_data_244_1 = mem_244_1_R0_data;
  wire [7:0] R0_data_244_2 = mem_244_2_R0_data;
  wire [7:0] R0_data_244_3 = mem_244_3_R0_data;
  wire [7:0] R0_data_244_4 = mem_244_4_R0_data;
  wire [7:0] R0_data_244_5 = mem_244_5_R0_data;
  wire [7:0] R0_data_244_6 = mem_244_6_R0_data;
  wire [7:0] R0_data_244_7 = mem_244_7_R0_data;
  wire [63:0] R0_data_244 = {R0_data_244_7,R0_data_244_6,R0_data_244_5,R0_data_244_4,R0_data_244_3,R0_data_244_2,
    R0_data_244_1,R0_data_244_0};
  wire [7:0] R0_data_245_0 = mem_245_0_R0_data;
  wire [7:0] R0_data_245_1 = mem_245_1_R0_data;
  wire [7:0] R0_data_245_2 = mem_245_2_R0_data;
  wire [7:0] R0_data_245_3 = mem_245_3_R0_data;
  wire [7:0] R0_data_245_4 = mem_245_4_R0_data;
  wire [7:0] R0_data_245_5 = mem_245_5_R0_data;
  wire [7:0] R0_data_245_6 = mem_245_6_R0_data;
  wire [7:0] R0_data_245_7 = mem_245_7_R0_data;
  wire [63:0] R0_data_245 = {R0_data_245_7,R0_data_245_6,R0_data_245_5,R0_data_245_4,R0_data_245_3,R0_data_245_2,
    R0_data_245_1,R0_data_245_0};
  wire [7:0] R0_data_246_0 = mem_246_0_R0_data;
  wire [7:0] R0_data_246_1 = mem_246_1_R0_data;
  wire [7:0] R0_data_246_2 = mem_246_2_R0_data;
  wire [7:0] R0_data_246_3 = mem_246_3_R0_data;
  wire [7:0] R0_data_246_4 = mem_246_4_R0_data;
  wire [7:0] R0_data_246_5 = mem_246_5_R0_data;
  wire [7:0] R0_data_246_6 = mem_246_6_R0_data;
  wire [7:0] R0_data_246_7 = mem_246_7_R0_data;
  wire [63:0] R0_data_246 = {R0_data_246_7,R0_data_246_6,R0_data_246_5,R0_data_246_4,R0_data_246_3,R0_data_246_2,
    R0_data_246_1,R0_data_246_0};
  wire [7:0] R0_data_247_0 = mem_247_0_R0_data;
  wire [7:0] R0_data_247_1 = mem_247_1_R0_data;
  wire [7:0] R0_data_247_2 = mem_247_2_R0_data;
  wire [7:0] R0_data_247_3 = mem_247_3_R0_data;
  wire [7:0] R0_data_247_4 = mem_247_4_R0_data;
  wire [7:0] R0_data_247_5 = mem_247_5_R0_data;
  wire [7:0] R0_data_247_6 = mem_247_6_R0_data;
  wire [7:0] R0_data_247_7 = mem_247_7_R0_data;
  wire [63:0] R0_data_247 = {R0_data_247_7,R0_data_247_6,R0_data_247_5,R0_data_247_4,R0_data_247_3,R0_data_247_2,
    R0_data_247_1,R0_data_247_0};
  wire [7:0] R0_data_248_0 = mem_248_0_R0_data;
  wire [7:0] R0_data_248_1 = mem_248_1_R0_data;
  wire [7:0] R0_data_248_2 = mem_248_2_R0_data;
  wire [7:0] R0_data_248_3 = mem_248_3_R0_data;
  wire [7:0] R0_data_248_4 = mem_248_4_R0_data;
  wire [7:0] R0_data_248_5 = mem_248_5_R0_data;
  wire [7:0] R0_data_248_6 = mem_248_6_R0_data;
  wire [7:0] R0_data_248_7 = mem_248_7_R0_data;
  wire [63:0] R0_data_248 = {R0_data_248_7,R0_data_248_6,R0_data_248_5,R0_data_248_4,R0_data_248_3,R0_data_248_2,
    R0_data_248_1,R0_data_248_0};
  wire [7:0] R0_data_249_0 = mem_249_0_R0_data;
  wire [7:0] R0_data_249_1 = mem_249_1_R0_data;
  wire [7:0] R0_data_249_2 = mem_249_2_R0_data;
  wire [7:0] R0_data_249_3 = mem_249_3_R0_data;
  wire [7:0] R0_data_249_4 = mem_249_4_R0_data;
  wire [7:0] R0_data_249_5 = mem_249_5_R0_data;
  wire [7:0] R0_data_249_6 = mem_249_6_R0_data;
  wire [7:0] R0_data_249_7 = mem_249_7_R0_data;
  wire [63:0] R0_data_249 = {R0_data_249_7,R0_data_249_6,R0_data_249_5,R0_data_249_4,R0_data_249_3,R0_data_249_2,
    R0_data_249_1,R0_data_249_0};
  wire [7:0] R0_data_250_0 = mem_250_0_R0_data;
  wire [7:0] R0_data_250_1 = mem_250_1_R0_data;
  wire [7:0] R0_data_250_2 = mem_250_2_R0_data;
  wire [7:0] R0_data_250_3 = mem_250_3_R0_data;
  wire [7:0] R0_data_250_4 = mem_250_4_R0_data;
  wire [7:0] R0_data_250_5 = mem_250_5_R0_data;
  wire [7:0] R0_data_250_6 = mem_250_6_R0_data;
  wire [7:0] R0_data_250_7 = mem_250_7_R0_data;
  wire [63:0] R0_data_250 = {R0_data_250_7,R0_data_250_6,R0_data_250_5,R0_data_250_4,R0_data_250_3,R0_data_250_2,
    R0_data_250_1,R0_data_250_0};
  wire [7:0] R0_data_251_0 = mem_251_0_R0_data;
  wire [7:0] R0_data_251_1 = mem_251_1_R0_data;
  wire [7:0] R0_data_251_2 = mem_251_2_R0_data;
  wire [7:0] R0_data_251_3 = mem_251_3_R0_data;
  wire [7:0] R0_data_251_4 = mem_251_4_R0_data;
  wire [7:0] R0_data_251_5 = mem_251_5_R0_data;
  wire [7:0] R0_data_251_6 = mem_251_6_R0_data;
  wire [7:0] R0_data_251_7 = mem_251_7_R0_data;
  wire [63:0] R0_data_251 = {R0_data_251_7,R0_data_251_6,R0_data_251_5,R0_data_251_4,R0_data_251_3,R0_data_251_2,
    R0_data_251_1,R0_data_251_0};
  wire [7:0] R0_data_252_0 = mem_252_0_R0_data;
  wire [7:0] R0_data_252_1 = mem_252_1_R0_data;
  wire [7:0] R0_data_252_2 = mem_252_2_R0_data;
  wire [7:0] R0_data_252_3 = mem_252_3_R0_data;
  wire [7:0] R0_data_252_4 = mem_252_4_R0_data;
  wire [7:0] R0_data_252_5 = mem_252_5_R0_data;
  wire [7:0] R0_data_252_6 = mem_252_6_R0_data;
  wire [7:0] R0_data_252_7 = mem_252_7_R0_data;
  wire [63:0] R0_data_252 = {R0_data_252_7,R0_data_252_6,R0_data_252_5,R0_data_252_4,R0_data_252_3,R0_data_252_2,
    R0_data_252_1,R0_data_252_0};
  wire [7:0] R0_data_253_0 = mem_253_0_R0_data;
  wire [7:0] R0_data_253_1 = mem_253_1_R0_data;
  wire [7:0] R0_data_253_2 = mem_253_2_R0_data;
  wire [7:0] R0_data_253_3 = mem_253_3_R0_data;
  wire [7:0] R0_data_253_4 = mem_253_4_R0_data;
  wire [7:0] R0_data_253_5 = mem_253_5_R0_data;
  wire [7:0] R0_data_253_6 = mem_253_6_R0_data;
  wire [7:0] R0_data_253_7 = mem_253_7_R0_data;
  wire [63:0] R0_data_253 = {R0_data_253_7,R0_data_253_6,R0_data_253_5,R0_data_253_4,R0_data_253_3,R0_data_253_2,
    R0_data_253_1,R0_data_253_0};
  wire [7:0] R0_data_254_0 = mem_254_0_R0_data;
  wire [7:0] R0_data_254_1 = mem_254_1_R0_data;
  wire [7:0] R0_data_254_2 = mem_254_2_R0_data;
  wire [7:0] R0_data_254_3 = mem_254_3_R0_data;
  wire [7:0] R0_data_254_4 = mem_254_4_R0_data;
  wire [7:0] R0_data_254_5 = mem_254_5_R0_data;
  wire [7:0] R0_data_254_6 = mem_254_6_R0_data;
  wire [7:0] R0_data_254_7 = mem_254_7_R0_data;
  wire [63:0] R0_data_254 = {R0_data_254_7,R0_data_254_6,R0_data_254_5,R0_data_254_4,R0_data_254_3,R0_data_254_2,
    R0_data_254_1,R0_data_254_0};
  wire [7:0] R0_data_255_0 = mem_255_0_R0_data;
  wire [7:0] R0_data_255_1 = mem_255_1_R0_data;
  wire [7:0] R0_data_255_2 = mem_255_2_R0_data;
  wire [7:0] R0_data_255_3 = mem_255_3_R0_data;
  wire [7:0] R0_data_255_4 = mem_255_4_R0_data;
  wire [7:0] R0_data_255_5 = mem_255_5_R0_data;
  wire [7:0] R0_data_255_6 = mem_255_6_R0_data;
  wire [7:0] R0_data_255_7 = mem_255_7_R0_data;
  wire [63:0] R0_data_255 = {R0_data_255_7,R0_data_255_6,R0_data_255_5,R0_data_255_4,R0_data_255_3,R0_data_255_2,
    R0_data_255_1,R0_data_255_0};
  split_mem_0_ext mem_0_0 (
    .R0_addr(mem_0_0_R0_addr),
    .R0_clk(mem_0_0_R0_clk),
    .R0_data(mem_0_0_R0_data),
    .R0_en(mem_0_0_R0_en),
    .W0_addr(mem_0_0_W0_addr),
    .W0_clk(mem_0_0_W0_clk),
    .W0_data(mem_0_0_W0_data),
    .W0_en(mem_0_0_W0_en),
    .W0_mask(mem_0_0_W0_mask)
  );
  split_mem_0_ext mem_0_1 (
    .R0_addr(mem_0_1_R0_addr),
    .R0_clk(mem_0_1_R0_clk),
    .R0_data(mem_0_1_R0_data),
    .R0_en(mem_0_1_R0_en),
    .W0_addr(mem_0_1_W0_addr),
    .W0_clk(mem_0_1_W0_clk),
    .W0_data(mem_0_1_W0_data),
    .W0_en(mem_0_1_W0_en),
    .W0_mask(mem_0_1_W0_mask)
  );
  split_mem_0_ext mem_0_2 (
    .R0_addr(mem_0_2_R0_addr),
    .R0_clk(mem_0_2_R0_clk),
    .R0_data(mem_0_2_R0_data),
    .R0_en(mem_0_2_R0_en),
    .W0_addr(mem_0_2_W0_addr),
    .W0_clk(mem_0_2_W0_clk),
    .W0_data(mem_0_2_W0_data),
    .W0_en(mem_0_2_W0_en),
    .W0_mask(mem_0_2_W0_mask)
  );
  split_mem_0_ext mem_0_3 (
    .R0_addr(mem_0_3_R0_addr),
    .R0_clk(mem_0_3_R0_clk),
    .R0_data(mem_0_3_R0_data),
    .R0_en(mem_0_3_R0_en),
    .W0_addr(mem_0_3_W0_addr),
    .W0_clk(mem_0_3_W0_clk),
    .W0_data(mem_0_3_W0_data),
    .W0_en(mem_0_3_W0_en),
    .W0_mask(mem_0_3_W0_mask)
  );
  split_mem_0_ext mem_0_4 (
    .R0_addr(mem_0_4_R0_addr),
    .R0_clk(mem_0_4_R0_clk),
    .R0_data(mem_0_4_R0_data),
    .R0_en(mem_0_4_R0_en),
    .W0_addr(mem_0_4_W0_addr),
    .W0_clk(mem_0_4_W0_clk),
    .W0_data(mem_0_4_W0_data),
    .W0_en(mem_0_4_W0_en),
    .W0_mask(mem_0_4_W0_mask)
  );
  split_mem_0_ext mem_0_5 (
    .R0_addr(mem_0_5_R0_addr),
    .R0_clk(mem_0_5_R0_clk),
    .R0_data(mem_0_5_R0_data),
    .R0_en(mem_0_5_R0_en),
    .W0_addr(mem_0_5_W0_addr),
    .W0_clk(mem_0_5_W0_clk),
    .W0_data(mem_0_5_W0_data),
    .W0_en(mem_0_5_W0_en),
    .W0_mask(mem_0_5_W0_mask)
  );
  split_mem_0_ext mem_0_6 (
    .R0_addr(mem_0_6_R0_addr),
    .R0_clk(mem_0_6_R0_clk),
    .R0_data(mem_0_6_R0_data),
    .R0_en(mem_0_6_R0_en),
    .W0_addr(mem_0_6_W0_addr),
    .W0_clk(mem_0_6_W0_clk),
    .W0_data(mem_0_6_W0_data),
    .W0_en(mem_0_6_W0_en),
    .W0_mask(mem_0_6_W0_mask)
  );
  split_mem_0_ext mem_0_7 (
    .R0_addr(mem_0_7_R0_addr),
    .R0_clk(mem_0_7_R0_clk),
    .R0_data(mem_0_7_R0_data),
    .R0_en(mem_0_7_R0_en),
    .W0_addr(mem_0_7_W0_addr),
    .W0_clk(mem_0_7_W0_clk),
    .W0_data(mem_0_7_W0_data),
    .W0_en(mem_0_7_W0_en),
    .W0_mask(mem_0_7_W0_mask)
  );
  split_mem_0_ext mem_1_0 (
    .R0_addr(mem_1_0_R0_addr),
    .R0_clk(mem_1_0_R0_clk),
    .R0_data(mem_1_0_R0_data),
    .R0_en(mem_1_0_R0_en),
    .W0_addr(mem_1_0_W0_addr),
    .W0_clk(mem_1_0_W0_clk),
    .W0_data(mem_1_0_W0_data),
    .W0_en(mem_1_0_W0_en),
    .W0_mask(mem_1_0_W0_mask)
  );
  split_mem_0_ext mem_1_1 (
    .R0_addr(mem_1_1_R0_addr),
    .R0_clk(mem_1_1_R0_clk),
    .R0_data(mem_1_1_R0_data),
    .R0_en(mem_1_1_R0_en),
    .W0_addr(mem_1_1_W0_addr),
    .W0_clk(mem_1_1_W0_clk),
    .W0_data(mem_1_1_W0_data),
    .W0_en(mem_1_1_W0_en),
    .W0_mask(mem_1_1_W0_mask)
  );
  split_mem_0_ext mem_1_2 (
    .R0_addr(mem_1_2_R0_addr),
    .R0_clk(mem_1_2_R0_clk),
    .R0_data(mem_1_2_R0_data),
    .R0_en(mem_1_2_R0_en),
    .W0_addr(mem_1_2_W0_addr),
    .W0_clk(mem_1_2_W0_clk),
    .W0_data(mem_1_2_W0_data),
    .W0_en(mem_1_2_W0_en),
    .W0_mask(mem_1_2_W0_mask)
  );
  split_mem_0_ext mem_1_3 (
    .R0_addr(mem_1_3_R0_addr),
    .R0_clk(mem_1_3_R0_clk),
    .R0_data(mem_1_3_R0_data),
    .R0_en(mem_1_3_R0_en),
    .W0_addr(mem_1_3_W0_addr),
    .W0_clk(mem_1_3_W0_clk),
    .W0_data(mem_1_3_W0_data),
    .W0_en(mem_1_3_W0_en),
    .W0_mask(mem_1_3_W0_mask)
  );
  split_mem_0_ext mem_1_4 (
    .R0_addr(mem_1_4_R0_addr),
    .R0_clk(mem_1_4_R0_clk),
    .R0_data(mem_1_4_R0_data),
    .R0_en(mem_1_4_R0_en),
    .W0_addr(mem_1_4_W0_addr),
    .W0_clk(mem_1_4_W0_clk),
    .W0_data(mem_1_4_W0_data),
    .W0_en(mem_1_4_W0_en),
    .W0_mask(mem_1_4_W0_mask)
  );
  split_mem_0_ext mem_1_5 (
    .R0_addr(mem_1_5_R0_addr),
    .R0_clk(mem_1_5_R0_clk),
    .R0_data(mem_1_5_R0_data),
    .R0_en(mem_1_5_R0_en),
    .W0_addr(mem_1_5_W0_addr),
    .W0_clk(mem_1_5_W0_clk),
    .W0_data(mem_1_5_W0_data),
    .W0_en(mem_1_5_W0_en),
    .W0_mask(mem_1_5_W0_mask)
  );
  split_mem_0_ext mem_1_6 (
    .R0_addr(mem_1_6_R0_addr),
    .R0_clk(mem_1_6_R0_clk),
    .R0_data(mem_1_6_R0_data),
    .R0_en(mem_1_6_R0_en),
    .W0_addr(mem_1_6_W0_addr),
    .W0_clk(mem_1_6_W0_clk),
    .W0_data(mem_1_6_W0_data),
    .W0_en(mem_1_6_W0_en),
    .W0_mask(mem_1_6_W0_mask)
  );
  split_mem_0_ext mem_1_7 (
    .R0_addr(mem_1_7_R0_addr),
    .R0_clk(mem_1_7_R0_clk),
    .R0_data(mem_1_7_R0_data),
    .R0_en(mem_1_7_R0_en),
    .W0_addr(mem_1_7_W0_addr),
    .W0_clk(mem_1_7_W0_clk),
    .W0_data(mem_1_7_W0_data),
    .W0_en(mem_1_7_W0_en),
    .W0_mask(mem_1_7_W0_mask)
  );
  split_mem_0_ext mem_2_0 (
    .R0_addr(mem_2_0_R0_addr),
    .R0_clk(mem_2_0_R0_clk),
    .R0_data(mem_2_0_R0_data),
    .R0_en(mem_2_0_R0_en),
    .W0_addr(mem_2_0_W0_addr),
    .W0_clk(mem_2_0_W0_clk),
    .W0_data(mem_2_0_W0_data),
    .W0_en(mem_2_0_W0_en),
    .W0_mask(mem_2_0_W0_mask)
  );
  split_mem_0_ext mem_2_1 (
    .R0_addr(mem_2_1_R0_addr),
    .R0_clk(mem_2_1_R0_clk),
    .R0_data(mem_2_1_R0_data),
    .R0_en(mem_2_1_R0_en),
    .W0_addr(mem_2_1_W0_addr),
    .W0_clk(mem_2_1_W0_clk),
    .W0_data(mem_2_1_W0_data),
    .W0_en(mem_2_1_W0_en),
    .W0_mask(mem_2_1_W0_mask)
  );
  split_mem_0_ext mem_2_2 (
    .R0_addr(mem_2_2_R0_addr),
    .R0_clk(mem_2_2_R0_clk),
    .R0_data(mem_2_2_R0_data),
    .R0_en(mem_2_2_R0_en),
    .W0_addr(mem_2_2_W0_addr),
    .W0_clk(mem_2_2_W0_clk),
    .W0_data(mem_2_2_W0_data),
    .W0_en(mem_2_2_W0_en),
    .W0_mask(mem_2_2_W0_mask)
  );
  split_mem_0_ext mem_2_3 (
    .R0_addr(mem_2_3_R0_addr),
    .R0_clk(mem_2_3_R0_clk),
    .R0_data(mem_2_3_R0_data),
    .R0_en(mem_2_3_R0_en),
    .W0_addr(mem_2_3_W0_addr),
    .W0_clk(mem_2_3_W0_clk),
    .W0_data(mem_2_3_W0_data),
    .W0_en(mem_2_3_W0_en),
    .W0_mask(mem_2_3_W0_mask)
  );
  split_mem_0_ext mem_2_4 (
    .R0_addr(mem_2_4_R0_addr),
    .R0_clk(mem_2_4_R0_clk),
    .R0_data(mem_2_4_R0_data),
    .R0_en(mem_2_4_R0_en),
    .W0_addr(mem_2_4_W0_addr),
    .W0_clk(mem_2_4_W0_clk),
    .W0_data(mem_2_4_W0_data),
    .W0_en(mem_2_4_W0_en),
    .W0_mask(mem_2_4_W0_mask)
  );
  split_mem_0_ext mem_2_5 (
    .R0_addr(mem_2_5_R0_addr),
    .R0_clk(mem_2_5_R0_clk),
    .R0_data(mem_2_5_R0_data),
    .R0_en(mem_2_5_R0_en),
    .W0_addr(mem_2_5_W0_addr),
    .W0_clk(mem_2_5_W0_clk),
    .W0_data(mem_2_5_W0_data),
    .W0_en(mem_2_5_W0_en),
    .W0_mask(mem_2_5_W0_mask)
  );
  split_mem_0_ext mem_2_6 (
    .R0_addr(mem_2_6_R0_addr),
    .R0_clk(mem_2_6_R0_clk),
    .R0_data(mem_2_6_R0_data),
    .R0_en(mem_2_6_R0_en),
    .W0_addr(mem_2_6_W0_addr),
    .W0_clk(mem_2_6_W0_clk),
    .W0_data(mem_2_6_W0_data),
    .W0_en(mem_2_6_W0_en),
    .W0_mask(mem_2_6_W0_mask)
  );
  split_mem_0_ext mem_2_7 (
    .R0_addr(mem_2_7_R0_addr),
    .R0_clk(mem_2_7_R0_clk),
    .R0_data(mem_2_7_R0_data),
    .R0_en(mem_2_7_R0_en),
    .W0_addr(mem_2_7_W0_addr),
    .W0_clk(mem_2_7_W0_clk),
    .W0_data(mem_2_7_W0_data),
    .W0_en(mem_2_7_W0_en),
    .W0_mask(mem_2_7_W0_mask)
  );
  split_mem_0_ext mem_3_0 (
    .R0_addr(mem_3_0_R0_addr),
    .R0_clk(mem_3_0_R0_clk),
    .R0_data(mem_3_0_R0_data),
    .R0_en(mem_3_0_R0_en),
    .W0_addr(mem_3_0_W0_addr),
    .W0_clk(mem_3_0_W0_clk),
    .W0_data(mem_3_0_W0_data),
    .W0_en(mem_3_0_W0_en),
    .W0_mask(mem_3_0_W0_mask)
  );
  split_mem_0_ext mem_3_1 (
    .R0_addr(mem_3_1_R0_addr),
    .R0_clk(mem_3_1_R0_clk),
    .R0_data(mem_3_1_R0_data),
    .R0_en(mem_3_1_R0_en),
    .W0_addr(mem_3_1_W0_addr),
    .W0_clk(mem_3_1_W0_clk),
    .W0_data(mem_3_1_W0_data),
    .W0_en(mem_3_1_W0_en),
    .W0_mask(mem_3_1_W0_mask)
  );
  split_mem_0_ext mem_3_2 (
    .R0_addr(mem_3_2_R0_addr),
    .R0_clk(mem_3_2_R0_clk),
    .R0_data(mem_3_2_R0_data),
    .R0_en(mem_3_2_R0_en),
    .W0_addr(mem_3_2_W0_addr),
    .W0_clk(mem_3_2_W0_clk),
    .W0_data(mem_3_2_W0_data),
    .W0_en(mem_3_2_W0_en),
    .W0_mask(mem_3_2_W0_mask)
  );
  split_mem_0_ext mem_3_3 (
    .R0_addr(mem_3_3_R0_addr),
    .R0_clk(mem_3_3_R0_clk),
    .R0_data(mem_3_3_R0_data),
    .R0_en(mem_3_3_R0_en),
    .W0_addr(mem_3_3_W0_addr),
    .W0_clk(mem_3_3_W0_clk),
    .W0_data(mem_3_3_W0_data),
    .W0_en(mem_3_3_W0_en),
    .W0_mask(mem_3_3_W0_mask)
  );
  split_mem_0_ext mem_3_4 (
    .R0_addr(mem_3_4_R0_addr),
    .R0_clk(mem_3_4_R0_clk),
    .R0_data(mem_3_4_R0_data),
    .R0_en(mem_3_4_R0_en),
    .W0_addr(mem_3_4_W0_addr),
    .W0_clk(mem_3_4_W0_clk),
    .W0_data(mem_3_4_W0_data),
    .W0_en(mem_3_4_W0_en),
    .W0_mask(mem_3_4_W0_mask)
  );
  split_mem_0_ext mem_3_5 (
    .R0_addr(mem_3_5_R0_addr),
    .R0_clk(mem_3_5_R0_clk),
    .R0_data(mem_3_5_R0_data),
    .R0_en(mem_3_5_R0_en),
    .W0_addr(mem_3_5_W0_addr),
    .W0_clk(mem_3_5_W0_clk),
    .W0_data(mem_3_5_W0_data),
    .W0_en(mem_3_5_W0_en),
    .W0_mask(mem_3_5_W0_mask)
  );
  split_mem_0_ext mem_3_6 (
    .R0_addr(mem_3_6_R0_addr),
    .R0_clk(mem_3_6_R0_clk),
    .R0_data(mem_3_6_R0_data),
    .R0_en(mem_3_6_R0_en),
    .W0_addr(mem_3_6_W0_addr),
    .W0_clk(mem_3_6_W0_clk),
    .W0_data(mem_3_6_W0_data),
    .W0_en(mem_3_6_W0_en),
    .W0_mask(mem_3_6_W0_mask)
  );
  split_mem_0_ext mem_3_7 (
    .R0_addr(mem_3_7_R0_addr),
    .R0_clk(mem_3_7_R0_clk),
    .R0_data(mem_3_7_R0_data),
    .R0_en(mem_3_7_R0_en),
    .W0_addr(mem_3_7_W0_addr),
    .W0_clk(mem_3_7_W0_clk),
    .W0_data(mem_3_7_W0_data),
    .W0_en(mem_3_7_W0_en),
    .W0_mask(mem_3_7_W0_mask)
  );
  split_mem_0_ext mem_4_0 (
    .R0_addr(mem_4_0_R0_addr),
    .R0_clk(mem_4_0_R0_clk),
    .R0_data(mem_4_0_R0_data),
    .R0_en(mem_4_0_R0_en),
    .W0_addr(mem_4_0_W0_addr),
    .W0_clk(mem_4_0_W0_clk),
    .W0_data(mem_4_0_W0_data),
    .W0_en(mem_4_0_W0_en),
    .W0_mask(mem_4_0_W0_mask)
  );
  split_mem_0_ext mem_4_1 (
    .R0_addr(mem_4_1_R0_addr),
    .R0_clk(mem_4_1_R0_clk),
    .R0_data(mem_4_1_R0_data),
    .R0_en(mem_4_1_R0_en),
    .W0_addr(mem_4_1_W0_addr),
    .W0_clk(mem_4_1_W0_clk),
    .W0_data(mem_4_1_W0_data),
    .W0_en(mem_4_1_W0_en),
    .W0_mask(mem_4_1_W0_mask)
  );
  split_mem_0_ext mem_4_2 (
    .R0_addr(mem_4_2_R0_addr),
    .R0_clk(mem_4_2_R0_clk),
    .R0_data(mem_4_2_R0_data),
    .R0_en(mem_4_2_R0_en),
    .W0_addr(mem_4_2_W0_addr),
    .W0_clk(mem_4_2_W0_clk),
    .W0_data(mem_4_2_W0_data),
    .W0_en(mem_4_2_W0_en),
    .W0_mask(mem_4_2_W0_mask)
  );
  split_mem_0_ext mem_4_3 (
    .R0_addr(mem_4_3_R0_addr),
    .R0_clk(mem_4_3_R0_clk),
    .R0_data(mem_4_3_R0_data),
    .R0_en(mem_4_3_R0_en),
    .W0_addr(mem_4_3_W0_addr),
    .W0_clk(mem_4_3_W0_clk),
    .W0_data(mem_4_3_W0_data),
    .W0_en(mem_4_3_W0_en),
    .W0_mask(mem_4_3_W0_mask)
  );
  split_mem_0_ext mem_4_4 (
    .R0_addr(mem_4_4_R0_addr),
    .R0_clk(mem_4_4_R0_clk),
    .R0_data(mem_4_4_R0_data),
    .R0_en(mem_4_4_R0_en),
    .W0_addr(mem_4_4_W0_addr),
    .W0_clk(mem_4_4_W0_clk),
    .W0_data(mem_4_4_W0_data),
    .W0_en(mem_4_4_W0_en),
    .W0_mask(mem_4_4_W0_mask)
  );
  split_mem_0_ext mem_4_5 (
    .R0_addr(mem_4_5_R0_addr),
    .R0_clk(mem_4_5_R0_clk),
    .R0_data(mem_4_5_R0_data),
    .R0_en(mem_4_5_R0_en),
    .W0_addr(mem_4_5_W0_addr),
    .W0_clk(mem_4_5_W0_clk),
    .W0_data(mem_4_5_W0_data),
    .W0_en(mem_4_5_W0_en),
    .W0_mask(mem_4_5_W0_mask)
  );
  split_mem_0_ext mem_4_6 (
    .R0_addr(mem_4_6_R0_addr),
    .R0_clk(mem_4_6_R0_clk),
    .R0_data(mem_4_6_R0_data),
    .R0_en(mem_4_6_R0_en),
    .W0_addr(mem_4_6_W0_addr),
    .W0_clk(mem_4_6_W0_clk),
    .W0_data(mem_4_6_W0_data),
    .W0_en(mem_4_6_W0_en),
    .W0_mask(mem_4_6_W0_mask)
  );
  split_mem_0_ext mem_4_7 (
    .R0_addr(mem_4_7_R0_addr),
    .R0_clk(mem_4_7_R0_clk),
    .R0_data(mem_4_7_R0_data),
    .R0_en(mem_4_7_R0_en),
    .W0_addr(mem_4_7_W0_addr),
    .W0_clk(mem_4_7_W0_clk),
    .W0_data(mem_4_7_W0_data),
    .W0_en(mem_4_7_W0_en),
    .W0_mask(mem_4_7_W0_mask)
  );
  split_mem_0_ext mem_5_0 (
    .R0_addr(mem_5_0_R0_addr),
    .R0_clk(mem_5_0_R0_clk),
    .R0_data(mem_5_0_R0_data),
    .R0_en(mem_5_0_R0_en),
    .W0_addr(mem_5_0_W0_addr),
    .W0_clk(mem_5_0_W0_clk),
    .W0_data(mem_5_0_W0_data),
    .W0_en(mem_5_0_W0_en),
    .W0_mask(mem_5_0_W0_mask)
  );
  split_mem_0_ext mem_5_1 (
    .R0_addr(mem_5_1_R0_addr),
    .R0_clk(mem_5_1_R0_clk),
    .R0_data(mem_5_1_R0_data),
    .R0_en(mem_5_1_R0_en),
    .W0_addr(mem_5_1_W0_addr),
    .W0_clk(mem_5_1_W0_clk),
    .W0_data(mem_5_1_W0_data),
    .W0_en(mem_5_1_W0_en),
    .W0_mask(mem_5_1_W0_mask)
  );
  split_mem_0_ext mem_5_2 (
    .R0_addr(mem_5_2_R0_addr),
    .R0_clk(mem_5_2_R0_clk),
    .R0_data(mem_5_2_R0_data),
    .R0_en(mem_5_2_R0_en),
    .W0_addr(mem_5_2_W0_addr),
    .W0_clk(mem_5_2_W0_clk),
    .W0_data(mem_5_2_W0_data),
    .W0_en(mem_5_2_W0_en),
    .W0_mask(mem_5_2_W0_mask)
  );
  split_mem_0_ext mem_5_3 (
    .R0_addr(mem_5_3_R0_addr),
    .R0_clk(mem_5_3_R0_clk),
    .R0_data(mem_5_3_R0_data),
    .R0_en(mem_5_3_R0_en),
    .W0_addr(mem_5_3_W0_addr),
    .W0_clk(mem_5_3_W0_clk),
    .W0_data(mem_5_3_W0_data),
    .W0_en(mem_5_3_W0_en),
    .W0_mask(mem_5_3_W0_mask)
  );
  split_mem_0_ext mem_5_4 (
    .R0_addr(mem_5_4_R0_addr),
    .R0_clk(mem_5_4_R0_clk),
    .R0_data(mem_5_4_R0_data),
    .R0_en(mem_5_4_R0_en),
    .W0_addr(mem_5_4_W0_addr),
    .W0_clk(mem_5_4_W0_clk),
    .W0_data(mem_5_4_W0_data),
    .W0_en(mem_5_4_W0_en),
    .W0_mask(mem_5_4_W0_mask)
  );
  split_mem_0_ext mem_5_5 (
    .R0_addr(mem_5_5_R0_addr),
    .R0_clk(mem_5_5_R0_clk),
    .R0_data(mem_5_5_R0_data),
    .R0_en(mem_5_5_R0_en),
    .W0_addr(mem_5_5_W0_addr),
    .W0_clk(mem_5_5_W0_clk),
    .W0_data(mem_5_5_W0_data),
    .W0_en(mem_5_5_W0_en),
    .W0_mask(mem_5_5_W0_mask)
  );
  split_mem_0_ext mem_5_6 (
    .R0_addr(mem_5_6_R0_addr),
    .R0_clk(mem_5_6_R0_clk),
    .R0_data(mem_5_6_R0_data),
    .R0_en(mem_5_6_R0_en),
    .W0_addr(mem_5_6_W0_addr),
    .W0_clk(mem_5_6_W0_clk),
    .W0_data(mem_5_6_W0_data),
    .W0_en(mem_5_6_W0_en),
    .W0_mask(mem_5_6_W0_mask)
  );
  split_mem_0_ext mem_5_7 (
    .R0_addr(mem_5_7_R0_addr),
    .R0_clk(mem_5_7_R0_clk),
    .R0_data(mem_5_7_R0_data),
    .R0_en(mem_5_7_R0_en),
    .W0_addr(mem_5_7_W0_addr),
    .W0_clk(mem_5_7_W0_clk),
    .W0_data(mem_5_7_W0_data),
    .W0_en(mem_5_7_W0_en),
    .W0_mask(mem_5_7_W0_mask)
  );
  split_mem_0_ext mem_6_0 (
    .R0_addr(mem_6_0_R0_addr),
    .R0_clk(mem_6_0_R0_clk),
    .R0_data(mem_6_0_R0_data),
    .R0_en(mem_6_0_R0_en),
    .W0_addr(mem_6_0_W0_addr),
    .W0_clk(mem_6_0_W0_clk),
    .W0_data(mem_6_0_W0_data),
    .W0_en(mem_6_0_W0_en),
    .W0_mask(mem_6_0_W0_mask)
  );
  split_mem_0_ext mem_6_1 (
    .R0_addr(mem_6_1_R0_addr),
    .R0_clk(mem_6_1_R0_clk),
    .R0_data(mem_6_1_R0_data),
    .R0_en(mem_6_1_R0_en),
    .W0_addr(mem_6_1_W0_addr),
    .W0_clk(mem_6_1_W0_clk),
    .W0_data(mem_6_1_W0_data),
    .W0_en(mem_6_1_W0_en),
    .W0_mask(mem_6_1_W0_mask)
  );
  split_mem_0_ext mem_6_2 (
    .R0_addr(mem_6_2_R0_addr),
    .R0_clk(mem_6_2_R0_clk),
    .R0_data(mem_6_2_R0_data),
    .R0_en(mem_6_2_R0_en),
    .W0_addr(mem_6_2_W0_addr),
    .W0_clk(mem_6_2_W0_clk),
    .W0_data(mem_6_2_W0_data),
    .W0_en(mem_6_2_W0_en),
    .W0_mask(mem_6_2_W0_mask)
  );
  split_mem_0_ext mem_6_3 (
    .R0_addr(mem_6_3_R0_addr),
    .R0_clk(mem_6_3_R0_clk),
    .R0_data(mem_6_3_R0_data),
    .R0_en(mem_6_3_R0_en),
    .W0_addr(mem_6_3_W0_addr),
    .W0_clk(mem_6_3_W0_clk),
    .W0_data(mem_6_3_W0_data),
    .W0_en(mem_6_3_W0_en),
    .W0_mask(mem_6_3_W0_mask)
  );
  split_mem_0_ext mem_6_4 (
    .R0_addr(mem_6_4_R0_addr),
    .R0_clk(mem_6_4_R0_clk),
    .R0_data(mem_6_4_R0_data),
    .R0_en(mem_6_4_R0_en),
    .W0_addr(mem_6_4_W0_addr),
    .W0_clk(mem_6_4_W0_clk),
    .W0_data(mem_6_4_W0_data),
    .W0_en(mem_6_4_W0_en),
    .W0_mask(mem_6_4_W0_mask)
  );
  split_mem_0_ext mem_6_5 (
    .R0_addr(mem_6_5_R0_addr),
    .R0_clk(mem_6_5_R0_clk),
    .R0_data(mem_6_5_R0_data),
    .R0_en(mem_6_5_R0_en),
    .W0_addr(mem_6_5_W0_addr),
    .W0_clk(mem_6_5_W0_clk),
    .W0_data(mem_6_5_W0_data),
    .W0_en(mem_6_5_W0_en),
    .W0_mask(mem_6_5_W0_mask)
  );
  split_mem_0_ext mem_6_6 (
    .R0_addr(mem_6_6_R0_addr),
    .R0_clk(mem_6_6_R0_clk),
    .R0_data(mem_6_6_R0_data),
    .R0_en(mem_6_6_R0_en),
    .W0_addr(mem_6_6_W0_addr),
    .W0_clk(mem_6_6_W0_clk),
    .W0_data(mem_6_6_W0_data),
    .W0_en(mem_6_6_W0_en),
    .W0_mask(mem_6_6_W0_mask)
  );
  split_mem_0_ext mem_6_7 (
    .R0_addr(mem_6_7_R0_addr),
    .R0_clk(mem_6_7_R0_clk),
    .R0_data(mem_6_7_R0_data),
    .R0_en(mem_6_7_R0_en),
    .W0_addr(mem_6_7_W0_addr),
    .W0_clk(mem_6_7_W0_clk),
    .W0_data(mem_6_7_W0_data),
    .W0_en(mem_6_7_W0_en),
    .W0_mask(mem_6_7_W0_mask)
  );
  split_mem_0_ext mem_7_0 (
    .R0_addr(mem_7_0_R0_addr),
    .R0_clk(mem_7_0_R0_clk),
    .R0_data(mem_7_0_R0_data),
    .R0_en(mem_7_0_R0_en),
    .W0_addr(mem_7_0_W0_addr),
    .W0_clk(mem_7_0_W0_clk),
    .W0_data(mem_7_0_W0_data),
    .W0_en(mem_7_0_W0_en),
    .W0_mask(mem_7_0_W0_mask)
  );
  split_mem_0_ext mem_7_1 (
    .R0_addr(mem_7_1_R0_addr),
    .R0_clk(mem_7_1_R0_clk),
    .R0_data(mem_7_1_R0_data),
    .R0_en(mem_7_1_R0_en),
    .W0_addr(mem_7_1_W0_addr),
    .W0_clk(mem_7_1_W0_clk),
    .W0_data(mem_7_1_W0_data),
    .W0_en(mem_7_1_W0_en),
    .W0_mask(mem_7_1_W0_mask)
  );
  split_mem_0_ext mem_7_2 (
    .R0_addr(mem_7_2_R0_addr),
    .R0_clk(mem_7_2_R0_clk),
    .R0_data(mem_7_2_R0_data),
    .R0_en(mem_7_2_R0_en),
    .W0_addr(mem_7_2_W0_addr),
    .W0_clk(mem_7_2_W0_clk),
    .W0_data(mem_7_2_W0_data),
    .W0_en(mem_7_2_W0_en),
    .W0_mask(mem_7_2_W0_mask)
  );
  split_mem_0_ext mem_7_3 (
    .R0_addr(mem_7_3_R0_addr),
    .R0_clk(mem_7_3_R0_clk),
    .R0_data(mem_7_3_R0_data),
    .R0_en(mem_7_3_R0_en),
    .W0_addr(mem_7_3_W0_addr),
    .W0_clk(mem_7_3_W0_clk),
    .W0_data(mem_7_3_W0_data),
    .W0_en(mem_7_3_W0_en),
    .W0_mask(mem_7_3_W0_mask)
  );
  split_mem_0_ext mem_7_4 (
    .R0_addr(mem_7_4_R0_addr),
    .R0_clk(mem_7_4_R0_clk),
    .R0_data(mem_7_4_R0_data),
    .R0_en(mem_7_4_R0_en),
    .W0_addr(mem_7_4_W0_addr),
    .W0_clk(mem_7_4_W0_clk),
    .W0_data(mem_7_4_W0_data),
    .W0_en(mem_7_4_W0_en),
    .W0_mask(mem_7_4_W0_mask)
  );
  split_mem_0_ext mem_7_5 (
    .R0_addr(mem_7_5_R0_addr),
    .R0_clk(mem_7_5_R0_clk),
    .R0_data(mem_7_5_R0_data),
    .R0_en(mem_7_5_R0_en),
    .W0_addr(mem_7_5_W0_addr),
    .W0_clk(mem_7_5_W0_clk),
    .W0_data(mem_7_5_W0_data),
    .W0_en(mem_7_5_W0_en),
    .W0_mask(mem_7_5_W0_mask)
  );
  split_mem_0_ext mem_7_6 (
    .R0_addr(mem_7_6_R0_addr),
    .R0_clk(mem_7_6_R0_clk),
    .R0_data(mem_7_6_R0_data),
    .R0_en(mem_7_6_R0_en),
    .W0_addr(mem_7_6_W0_addr),
    .W0_clk(mem_7_6_W0_clk),
    .W0_data(mem_7_6_W0_data),
    .W0_en(mem_7_6_W0_en),
    .W0_mask(mem_7_6_W0_mask)
  );
  split_mem_0_ext mem_7_7 (
    .R0_addr(mem_7_7_R0_addr),
    .R0_clk(mem_7_7_R0_clk),
    .R0_data(mem_7_7_R0_data),
    .R0_en(mem_7_7_R0_en),
    .W0_addr(mem_7_7_W0_addr),
    .W0_clk(mem_7_7_W0_clk),
    .W0_data(mem_7_7_W0_data),
    .W0_en(mem_7_7_W0_en),
    .W0_mask(mem_7_7_W0_mask)
  );
  split_mem_0_ext mem_8_0 (
    .R0_addr(mem_8_0_R0_addr),
    .R0_clk(mem_8_0_R0_clk),
    .R0_data(mem_8_0_R0_data),
    .R0_en(mem_8_0_R0_en),
    .W0_addr(mem_8_0_W0_addr),
    .W0_clk(mem_8_0_W0_clk),
    .W0_data(mem_8_0_W0_data),
    .W0_en(mem_8_0_W0_en),
    .W0_mask(mem_8_0_W0_mask)
  );
  split_mem_0_ext mem_8_1 (
    .R0_addr(mem_8_1_R0_addr),
    .R0_clk(mem_8_1_R0_clk),
    .R0_data(mem_8_1_R0_data),
    .R0_en(mem_8_1_R0_en),
    .W0_addr(mem_8_1_W0_addr),
    .W0_clk(mem_8_1_W0_clk),
    .W0_data(mem_8_1_W0_data),
    .W0_en(mem_8_1_W0_en),
    .W0_mask(mem_8_1_W0_mask)
  );
  split_mem_0_ext mem_8_2 (
    .R0_addr(mem_8_2_R0_addr),
    .R0_clk(mem_8_2_R0_clk),
    .R0_data(mem_8_2_R0_data),
    .R0_en(mem_8_2_R0_en),
    .W0_addr(mem_8_2_W0_addr),
    .W0_clk(mem_8_2_W0_clk),
    .W0_data(mem_8_2_W0_data),
    .W0_en(mem_8_2_W0_en),
    .W0_mask(mem_8_2_W0_mask)
  );
  split_mem_0_ext mem_8_3 (
    .R0_addr(mem_8_3_R0_addr),
    .R0_clk(mem_8_3_R0_clk),
    .R0_data(mem_8_3_R0_data),
    .R0_en(mem_8_3_R0_en),
    .W0_addr(mem_8_3_W0_addr),
    .W0_clk(mem_8_3_W0_clk),
    .W0_data(mem_8_3_W0_data),
    .W0_en(mem_8_3_W0_en),
    .W0_mask(mem_8_3_W0_mask)
  );
  split_mem_0_ext mem_8_4 (
    .R0_addr(mem_8_4_R0_addr),
    .R0_clk(mem_8_4_R0_clk),
    .R0_data(mem_8_4_R0_data),
    .R0_en(mem_8_4_R0_en),
    .W0_addr(mem_8_4_W0_addr),
    .W0_clk(mem_8_4_W0_clk),
    .W0_data(mem_8_4_W0_data),
    .W0_en(mem_8_4_W0_en),
    .W0_mask(mem_8_4_W0_mask)
  );
  split_mem_0_ext mem_8_5 (
    .R0_addr(mem_8_5_R0_addr),
    .R0_clk(mem_8_5_R0_clk),
    .R0_data(mem_8_5_R0_data),
    .R0_en(mem_8_5_R0_en),
    .W0_addr(mem_8_5_W0_addr),
    .W0_clk(mem_8_5_W0_clk),
    .W0_data(mem_8_5_W0_data),
    .W0_en(mem_8_5_W0_en),
    .W0_mask(mem_8_5_W0_mask)
  );
  split_mem_0_ext mem_8_6 (
    .R0_addr(mem_8_6_R0_addr),
    .R0_clk(mem_8_6_R0_clk),
    .R0_data(mem_8_6_R0_data),
    .R0_en(mem_8_6_R0_en),
    .W0_addr(mem_8_6_W0_addr),
    .W0_clk(mem_8_6_W0_clk),
    .W0_data(mem_8_6_W0_data),
    .W0_en(mem_8_6_W0_en),
    .W0_mask(mem_8_6_W0_mask)
  );
  split_mem_0_ext mem_8_7 (
    .R0_addr(mem_8_7_R0_addr),
    .R0_clk(mem_8_7_R0_clk),
    .R0_data(mem_8_7_R0_data),
    .R0_en(mem_8_7_R0_en),
    .W0_addr(mem_8_7_W0_addr),
    .W0_clk(mem_8_7_W0_clk),
    .W0_data(mem_8_7_W0_data),
    .W0_en(mem_8_7_W0_en),
    .W0_mask(mem_8_7_W0_mask)
  );
  split_mem_0_ext mem_9_0 (
    .R0_addr(mem_9_0_R0_addr),
    .R0_clk(mem_9_0_R0_clk),
    .R0_data(mem_9_0_R0_data),
    .R0_en(mem_9_0_R0_en),
    .W0_addr(mem_9_0_W0_addr),
    .W0_clk(mem_9_0_W0_clk),
    .W0_data(mem_9_0_W0_data),
    .W0_en(mem_9_0_W0_en),
    .W0_mask(mem_9_0_W0_mask)
  );
  split_mem_0_ext mem_9_1 (
    .R0_addr(mem_9_1_R0_addr),
    .R0_clk(mem_9_1_R0_clk),
    .R0_data(mem_9_1_R0_data),
    .R0_en(mem_9_1_R0_en),
    .W0_addr(mem_9_1_W0_addr),
    .W0_clk(mem_9_1_W0_clk),
    .W0_data(mem_9_1_W0_data),
    .W0_en(mem_9_1_W0_en),
    .W0_mask(mem_9_1_W0_mask)
  );
  split_mem_0_ext mem_9_2 (
    .R0_addr(mem_9_2_R0_addr),
    .R0_clk(mem_9_2_R0_clk),
    .R0_data(mem_9_2_R0_data),
    .R0_en(mem_9_2_R0_en),
    .W0_addr(mem_9_2_W0_addr),
    .W0_clk(mem_9_2_W0_clk),
    .W0_data(mem_9_2_W0_data),
    .W0_en(mem_9_2_W0_en),
    .W0_mask(mem_9_2_W0_mask)
  );
  split_mem_0_ext mem_9_3 (
    .R0_addr(mem_9_3_R0_addr),
    .R0_clk(mem_9_3_R0_clk),
    .R0_data(mem_9_3_R0_data),
    .R0_en(mem_9_3_R0_en),
    .W0_addr(mem_9_3_W0_addr),
    .W0_clk(mem_9_3_W0_clk),
    .W0_data(mem_9_3_W0_data),
    .W0_en(mem_9_3_W0_en),
    .W0_mask(mem_9_3_W0_mask)
  );
  split_mem_0_ext mem_9_4 (
    .R0_addr(mem_9_4_R0_addr),
    .R0_clk(mem_9_4_R0_clk),
    .R0_data(mem_9_4_R0_data),
    .R0_en(mem_9_4_R0_en),
    .W0_addr(mem_9_4_W0_addr),
    .W0_clk(mem_9_4_W0_clk),
    .W0_data(mem_9_4_W0_data),
    .W0_en(mem_9_4_W0_en),
    .W0_mask(mem_9_4_W0_mask)
  );
  split_mem_0_ext mem_9_5 (
    .R0_addr(mem_9_5_R0_addr),
    .R0_clk(mem_9_5_R0_clk),
    .R0_data(mem_9_5_R0_data),
    .R0_en(mem_9_5_R0_en),
    .W0_addr(mem_9_5_W0_addr),
    .W0_clk(mem_9_5_W0_clk),
    .W0_data(mem_9_5_W0_data),
    .W0_en(mem_9_5_W0_en),
    .W0_mask(mem_9_5_W0_mask)
  );
  split_mem_0_ext mem_9_6 (
    .R0_addr(mem_9_6_R0_addr),
    .R0_clk(mem_9_6_R0_clk),
    .R0_data(mem_9_6_R0_data),
    .R0_en(mem_9_6_R0_en),
    .W0_addr(mem_9_6_W0_addr),
    .W0_clk(mem_9_6_W0_clk),
    .W0_data(mem_9_6_W0_data),
    .W0_en(mem_9_6_W0_en),
    .W0_mask(mem_9_6_W0_mask)
  );
  split_mem_0_ext mem_9_7 (
    .R0_addr(mem_9_7_R0_addr),
    .R0_clk(mem_9_7_R0_clk),
    .R0_data(mem_9_7_R0_data),
    .R0_en(mem_9_7_R0_en),
    .W0_addr(mem_9_7_W0_addr),
    .W0_clk(mem_9_7_W0_clk),
    .W0_data(mem_9_7_W0_data),
    .W0_en(mem_9_7_W0_en),
    .W0_mask(mem_9_7_W0_mask)
  );
  split_mem_0_ext mem_10_0 (
    .R0_addr(mem_10_0_R0_addr),
    .R0_clk(mem_10_0_R0_clk),
    .R0_data(mem_10_0_R0_data),
    .R0_en(mem_10_0_R0_en),
    .W0_addr(mem_10_0_W0_addr),
    .W0_clk(mem_10_0_W0_clk),
    .W0_data(mem_10_0_W0_data),
    .W0_en(mem_10_0_W0_en),
    .W0_mask(mem_10_0_W0_mask)
  );
  split_mem_0_ext mem_10_1 (
    .R0_addr(mem_10_1_R0_addr),
    .R0_clk(mem_10_1_R0_clk),
    .R0_data(mem_10_1_R0_data),
    .R0_en(mem_10_1_R0_en),
    .W0_addr(mem_10_1_W0_addr),
    .W0_clk(mem_10_1_W0_clk),
    .W0_data(mem_10_1_W0_data),
    .W0_en(mem_10_1_W0_en),
    .W0_mask(mem_10_1_W0_mask)
  );
  split_mem_0_ext mem_10_2 (
    .R0_addr(mem_10_2_R0_addr),
    .R0_clk(mem_10_2_R0_clk),
    .R0_data(mem_10_2_R0_data),
    .R0_en(mem_10_2_R0_en),
    .W0_addr(mem_10_2_W0_addr),
    .W0_clk(mem_10_2_W0_clk),
    .W0_data(mem_10_2_W0_data),
    .W0_en(mem_10_2_W0_en),
    .W0_mask(mem_10_2_W0_mask)
  );
  split_mem_0_ext mem_10_3 (
    .R0_addr(mem_10_3_R0_addr),
    .R0_clk(mem_10_3_R0_clk),
    .R0_data(mem_10_3_R0_data),
    .R0_en(mem_10_3_R0_en),
    .W0_addr(mem_10_3_W0_addr),
    .W0_clk(mem_10_3_W0_clk),
    .W0_data(mem_10_3_W0_data),
    .W0_en(mem_10_3_W0_en),
    .W0_mask(mem_10_3_W0_mask)
  );
  split_mem_0_ext mem_10_4 (
    .R0_addr(mem_10_4_R0_addr),
    .R0_clk(mem_10_4_R0_clk),
    .R0_data(mem_10_4_R0_data),
    .R0_en(mem_10_4_R0_en),
    .W0_addr(mem_10_4_W0_addr),
    .W0_clk(mem_10_4_W0_clk),
    .W0_data(mem_10_4_W0_data),
    .W0_en(mem_10_4_W0_en),
    .W0_mask(mem_10_4_W0_mask)
  );
  split_mem_0_ext mem_10_5 (
    .R0_addr(mem_10_5_R0_addr),
    .R0_clk(mem_10_5_R0_clk),
    .R0_data(mem_10_5_R0_data),
    .R0_en(mem_10_5_R0_en),
    .W0_addr(mem_10_5_W0_addr),
    .W0_clk(mem_10_5_W0_clk),
    .W0_data(mem_10_5_W0_data),
    .W0_en(mem_10_5_W0_en),
    .W0_mask(mem_10_5_W0_mask)
  );
  split_mem_0_ext mem_10_6 (
    .R0_addr(mem_10_6_R0_addr),
    .R0_clk(mem_10_6_R0_clk),
    .R0_data(mem_10_6_R0_data),
    .R0_en(mem_10_6_R0_en),
    .W0_addr(mem_10_6_W0_addr),
    .W0_clk(mem_10_6_W0_clk),
    .W0_data(mem_10_6_W0_data),
    .W0_en(mem_10_6_W0_en),
    .W0_mask(mem_10_6_W0_mask)
  );
  split_mem_0_ext mem_10_7 (
    .R0_addr(mem_10_7_R0_addr),
    .R0_clk(mem_10_7_R0_clk),
    .R0_data(mem_10_7_R0_data),
    .R0_en(mem_10_7_R0_en),
    .W0_addr(mem_10_7_W0_addr),
    .W0_clk(mem_10_7_W0_clk),
    .W0_data(mem_10_7_W0_data),
    .W0_en(mem_10_7_W0_en),
    .W0_mask(mem_10_7_W0_mask)
  );
  split_mem_0_ext mem_11_0 (
    .R0_addr(mem_11_0_R0_addr),
    .R0_clk(mem_11_0_R0_clk),
    .R0_data(mem_11_0_R0_data),
    .R0_en(mem_11_0_R0_en),
    .W0_addr(mem_11_0_W0_addr),
    .W0_clk(mem_11_0_W0_clk),
    .W0_data(mem_11_0_W0_data),
    .W0_en(mem_11_0_W0_en),
    .W0_mask(mem_11_0_W0_mask)
  );
  split_mem_0_ext mem_11_1 (
    .R0_addr(mem_11_1_R0_addr),
    .R0_clk(mem_11_1_R0_clk),
    .R0_data(mem_11_1_R0_data),
    .R0_en(mem_11_1_R0_en),
    .W0_addr(mem_11_1_W0_addr),
    .W0_clk(mem_11_1_W0_clk),
    .W0_data(mem_11_1_W0_data),
    .W0_en(mem_11_1_W0_en),
    .W0_mask(mem_11_1_W0_mask)
  );
  split_mem_0_ext mem_11_2 (
    .R0_addr(mem_11_2_R0_addr),
    .R0_clk(mem_11_2_R0_clk),
    .R0_data(mem_11_2_R0_data),
    .R0_en(mem_11_2_R0_en),
    .W0_addr(mem_11_2_W0_addr),
    .W0_clk(mem_11_2_W0_clk),
    .W0_data(mem_11_2_W0_data),
    .W0_en(mem_11_2_W0_en),
    .W0_mask(mem_11_2_W0_mask)
  );
  split_mem_0_ext mem_11_3 (
    .R0_addr(mem_11_3_R0_addr),
    .R0_clk(mem_11_3_R0_clk),
    .R0_data(mem_11_3_R0_data),
    .R0_en(mem_11_3_R0_en),
    .W0_addr(mem_11_3_W0_addr),
    .W0_clk(mem_11_3_W0_clk),
    .W0_data(mem_11_3_W0_data),
    .W0_en(mem_11_3_W0_en),
    .W0_mask(mem_11_3_W0_mask)
  );
  split_mem_0_ext mem_11_4 (
    .R0_addr(mem_11_4_R0_addr),
    .R0_clk(mem_11_4_R0_clk),
    .R0_data(mem_11_4_R0_data),
    .R0_en(mem_11_4_R0_en),
    .W0_addr(mem_11_4_W0_addr),
    .W0_clk(mem_11_4_W0_clk),
    .W0_data(mem_11_4_W0_data),
    .W0_en(mem_11_4_W0_en),
    .W0_mask(mem_11_4_W0_mask)
  );
  split_mem_0_ext mem_11_5 (
    .R0_addr(mem_11_5_R0_addr),
    .R0_clk(mem_11_5_R0_clk),
    .R0_data(mem_11_5_R0_data),
    .R0_en(mem_11_5_R0_en),
    .W0_addr(mem_11_5_W0_addr),
    .W0_clk(mem_11_5_W0_clk),
    .W0_data(mem_11_5_W0_data),
    .W0_en(mem_11_5_W0_en),
    .W0_mask(mem_11_5_W0_mask)
  );
  split_mem_0_ext mem_11_6 (
    .R0_addr(mem_11_6_R0_addr),
    .R0_clk(mem_11_6_R0_clk),
    .R0_data(mem_11_6_R0_data),
    .R0_en(mem_11_6_R0_en),
    .W0_addr(mem_11_6_W0_addr),
    .W0_clk(mem_11_6_W0_clk),
    .W0_data(mem_11_6_W0_data),
    .W0_en(mem_11_6_W0_en),
    .W0_mask(mem_11_6_W0_mask)
  );
  split_mem_0_ext mem_11_7 (
    .R0_addr(mem_11_7_R0_addr),
    .R0_clk(mem_11_7_R0_clk),
    .R0_data(mem_11_7_R0_data),
    .R0_en(mem_11_7_R0_en),
    .W0_addr(mem_11_7_W0_addr),
    .W0_clk(mem_11_7_W0_clk),
    .W0_data(mem_11_7_W0_data),
    .W0_en(mem_11_7_W0_en),
    .W0_mask(mem_11_7_W0_mask)
  );
  split_mem_0_ext mem_12_0 (
    .R0_addr(mem_12_0_R0_addr),
    .R0_clk(mem_12_0_R0_clk),
    .R0_data(mem_12_0_R0_data),
    .R0_en(mem_12_0_R0_en),
    .W0_addr(mem_12_0_W0_addr),
    .W0_clk(mem_12_0_W0_clk),
    .W0_data(mem_12_0_W0_data),
    .W0_en(mem_12_0_W0_en),
    .W0_mask(mem_12_0_W0_mask)
  );
  split_mem_0_ext mem_12_1 (
    .R0_addr(mem_12_1_R0_addr),
    .R0_clk(mem_12_1_R0_clk),
    .R0_data(mem_12_1_R0_data),
    .R0_en(mem_12_1_R0_en),
    .W0_addr(mem_12_1_W0_addr),
    .W0_clk(mem_12_1_W0_clk),
    .W0_data(mem_12_1_W0_data),
    .W0_en(mem_12_1_W0_en),
    .W0_mask(mem_12_1_W0_mask)
  );
  split_mem_0_ext mem_12_2 (
    .R0_addr(mem_12_2_R0_addr),
    .R0_clk(mem_12_2_R0_clk),
    .R0_data(mem_12_2_R0_data),
    .R0_en(mem_12_2_R0_en),
    .W0_addr(mem_12_2_W0_addr),
    .W0_clk(mem_12_2_W0_clk),
    .W0_data(mem_12_2_W0_data),
    .W0_en(mem_12_2_W0_en),
    .W0_mask(mem_12_2_W0_mask)
  );
  split_mem_0_ext mem_12_3 (
    .R0_addr(mem_12_3_R0_addr),
    .R0_clk(mem_12_3_R0_clk),
    .R0_data(mem_12_3_R0_data),
    .R0_en(mem_12_3_R0_en),
    .W0_addr(mem_12_3_W0_addr),
    .W0_clk(mem_12_3_W0_clk),
    .W0_data(mem_12_3_W0_data),
    .W0_en(mem_12_3_W0_en),
    .W0_mask(mem_12_3_W0_mask)
  );
  split_mem_0_ext mem_12_4 (
    .R0_addr(mem_12_4_R0_addr),
    .R0_clk(mem_12_4_R0_clk),
    .R0_data(mem_12_4_R0_data),
    .R0_en(mem_12_4_R0_en),
    .W0_addr(mem_12_4_W0_addr),
    .W0_clk(mem_12_4_W0_clk),
    .W0_data(mem_12_4_W0_data),
    .W0_en(mem_12_4_W0_en),
    .W0_mask(mem_12_4_W0_mask)
  );
  split_mem_0_ext mem_12_5 (
    .R0_addr(mem_12_5_R0_addr),
    .R0_clk(mem_12_5_R0_clk),
    .R0_data(mem_12_5_R0_data),
    .R0_en(mem_12_5_R0_en),
    .W0_addr(mem_12_5_W0_addr),
    .W0_clk(mem_12_5_W0_clk),
    .W0_data(mem_12_5_W0_data),
    .W0_en(mem_12_5_W0_en),
    .W0_mask(mem_12_5_W0_mask)
  );
  split_mem_0_ext mem_12_6 (
    .R0_addr(mem_12_6_R0_addr),
    .R0_clk(mem_12_6_R0_clk),
    .R0_data(mem_12_6_R0_data),
    .R0_en(mem_12_6_R0_en),
    .W0_addr(mem_12_6_W0_addr),
    .W0_clk(mem_12_6_W0_clk),
    .W0_data(mem_12_6_W0_data),
    .W0_en(mem_12_6_W0_en),
    .W0_mask(mem_12_6_W0_mask)
  );
  split_mem_0_ext mem_12_7 (
    .R0_addr(mem_12_7_R0_addr),
    .R0_clk(mem_12_7_R0_clk),
    .R0_data(mem_12_7_R0_data),
    .R0_en(mem_12_7_R0_en),
    .W0_addr(mem_12_7_W0_addr),
    .W0_clk(mem_12_7_W0_clk),
    .W0_data(mem_12_7_W0_data),
    .W0_en(mem_12_7_W0_en),
    .W0_mask(mem_12_7_W0_mask)
  );
  split_mem_0_ext mem_13_0 (
    .R0_addr(mem_13_0_R0_addr),
    .R0_clk(mem_13_0_R0_clk),
    .R0_data(mem_13_0_R0_data),
    .R0_en(mem_13_0_R0_en),
    .W0_addr(mem_13_0_W0_addr),
    .W0_clk(mem_13_0_W0_clk),
    .W0_data(mem_13_0_W0_data),
    .W0_en(mem_13_0_W0_en),
    .W0_mask(mem_13_0_W0_mask)
  );
  split_mem_0_ext mem_13_1 (
    .R0_addr(mem_13_1_R0_addr),
    .R0_clk(mem_13_1_R0_clk),
    .R0_data(mem_13_1_R0_data),
    .R0_en(mem_13_1_R0_en),
    .W0_addr(mem_13_1_W0_addr),
    .W0_clk(mem_13_1_W0_clk),
    .W0_data(mem_13_1_W0_data),
    .W0_en(mem_13_1_W0_en),
    .W0_mask(mem_13_1_W0_mask)
  );
  split_mem_0_ext mem_13_2 (
    .R0_addr(mem_13_2_R0_addr),
    .R0_clk(mem_13_2_R0_clk),
    .R0_data(mem_13_2_R0_data),
    .R0_en(mem_13_2_R0_en),
    .W0_addr(mem_13_2_W0_addr),
    .W0_clk(mem_13_2_W0_clk),
    .W0_data(mem_13_2_W0_data),
    .W0_en(mem_13_2_W0_en),
    .W0_mask(mem_13_2_W0_mask)
  );
  split_mem_0_ext mem_13_3 (
    .R0_addr(mem_13_3_R0_addr),
    .R0_clk(mem_13_3_R0_clk),
    .R0_data(mem_13_3_R0_data),
    .R0_en(mem_13_3_R0_en),
    .W0_addr(mem_13_3_W0_addr),
    .W0_clk(mem_13_3_W0_clk),
    .W0_data(mem_13_3_W0_data),
    .W0_en(mem_13_3_W0_en),
    .W0_mask(mem_13_3_W0_mask)
  );
  split_mem_0_ext mem_13_4 (
    .R0_addr(mem_13_4_R0_addr),
    .R0_clk(mem_13_4_R0_clk),
    .R0_data(mem_13_4_R0_data),
    .R0_en(mem_13_4_R0_en),
    .W0_addr(mem_13_4_W0_addr),
    .W0_clk(mem_13_4_W0_clk),
    .W0_data(mem_13_4_W0_data),
    .W0_en(mem_13_4_W0_en),
    .W0_mask(mem_13_4_W0_mask)
  );
  split_mem_0_ext mem_13_5 (
    .R0_addr(mem_13_5_R0_addr),
    .R0_clk(mem_13_5_R0_clk),
    .R0_data(mem_13_5_R0_data),
    .R0_en(mem_13_5_R0_en),
    .W0_addr(mem_13_5_W0_addr),
    .W0_clk(mem_13_5_W0_clk),
    .W0_data(mem_13_5_W0_data),
    .W0_en(mem_13_5_W0_en),
    .W0_mask(mem_13_5_W0_mask)
  );
  split_mem_0_ext mem_13_6 (
    .R0_addr(mem_13_6_R0_addr),
    .R0_clk(mem_13_6_R0_clk),
    .R0_data(mem_13_6_R0_data),
    .R0_en(mem_13_6_R0_en),
    .W0_addr(mem_13_6_W0_addr),
    .W0_clk(mem_13_6_W0_clk),
    .W0_data(mem_13_6_W0_data),
    .W0_en(mem_13_6_W0_en),
    .W0_mask(mem_13_6_W0_mask)
  );
  split_mem_0_ext mem_13_7 (
    .R0_addr(mem_13_7_R0_addr),
    .R0_clk(mem_13_7_R0_clk),
    .R0_data(mem_13_7_R0_data),
    .R0_en(mem_13_7_R0_en),
    .W0_addr(mem_13_7_W0_addr),
    .W0_clk(mem_13_7_W0_clk),
    .W0_data(mem_13_7_W0_data),
    .W0_en(mem_13_7_W0_en),
    .W0_mask(mem_13_7_W0_mask)
  );
  split_mem_0_ext mem_14_0 (
    .R0_addr(mem_14_0_R0_addr),
    .R0_clk(mem_14_0_R0_clk),
    .R0_data(mem_14_0_R0_data),
    .R0_en(mem_14_0_R0_en),
    .W0_addr(mem_14_0_W0_addr),
    .W0_clk(mem_14_0_W0_clk),
    .W0_data(mem_14_0_W0_data),
    .W0_en(mem_14_0_W0_en),
    .W0_mask(mem_14_0_W0_mask)
  );
  split_mem_0_ext mem_14_1 (
    .R0_addr(mem_14_1_R0_addr),
    .R0_clk(mem_14_1_R0_clk),
    .R0_data(mem_14_1_R0_data),
    .R0_en(mem_14_1_R0_en),
    .W0_addr(mem_14_1_W0_addr),
    .W0_clk(mem_14_1_W0_clk),
    .W0_data(mem_14_1_W0_data),
    .W0_en(mem_14_1_W0_en),
    .W0_mask(mem_14_1_W0_mask)
  );
  split_mem_0_ext mem_14_2 (
    .R0_addr(mem_14_2_R0_addr),
    .R0_clk(mem_14_2_R0_clk),
    .R0_data(mem_14_2_R0_data),
    .R0_en(mem_14_2_R0_en),
    .W0_addr(mem_14_2_W0_addr),
    .W0_clk(mem_14_2_W0_clk),
    .W0_data(mem_14_2_W0_data),
    .W0_en(mem_14_2_W0_en),
    .W0_mask(mem_14_2_W0_mask)
  );
  split_mem_0_ext mem_14_3 (
    .R0_addr(mem_14_3_R0_addr),
    .R0_clk(mem_14_3_R0_clk),
    .R0_data(mem_14_3_R0_data),
    .R0_en(mem_14_3_R0_en),
    .W0_addr(mem_14_3_W0_addr),
    .W0_clk(mem_14_3_W0_clk),
    .W0_data(mem_14_3_W0_data),
    .W0_en(mem_14_3_W0_en),
    .W0_mask(mem_14_3_W0_mask)
  );
  split_mem_0_ext mem_14_4 (
    .R0_addr(mem_14_4_R0_addr),
    .R0_clk(mem_14_4_R0_clk),
    .R0_data(mem_14_4_R0_data),
    .R0_en(mem_14_4_R0_en),
    .W0_addr(mem_14_4_W0_addr),
    .W0_clk(mem_14_4_W0_clk),
    .W0_data(mem_14_4_W0_data),
    .W0_en(mem_14_4_W0_en),
    .W0_mask(mem_14_4_W0_mask)
  );
  split_mem_0_ext mem_14_5 (
    .R0_addr(mem_14_5_R0_addr),
    .R0_clk(mem_14_5_R0_clk),
    .R0_data(mem_14_5_R0_data),
    .R0_en(mem_14_5_R0_en),
    .W0_addr(mem_14_5_W0_addr),
    .W0_clk(mem_14_5_W0_clk),
    .W0_data(mem_14_5_W0_data),
    .W0_en(mem_14_5_W0_en),
    .W0_mask(mem_14_5_W0_mask)
  );
  split_mem_0_ext mem_14_6 (
    .R0_addr(mem_14_6_R0_addr),
    .R0_clk(mem_14_6_R0_clk),
    .R0_data(mem_14_6_R0_data),
    .R0_en(mem_14_6_R0_en),
    .W0_addr(mem_14_6_W0_addr),
    .W0_clk(mem_14_6_W0_clk),
    .W0_data(mem_14_6_W0_data),
    .W0_en(mem_14_6_W0_en),
    .W0_mask(mem_14_6_W0_mask)
  );
  split_mem_0_ext mem_14_7 (
    .R0_addr(mem_14_7_R0_addr),
    .R0_clk(mem_14_7_R0_clk),
    .R0_data(mem_14_7_R0_data),
    .R0_en(mem_14_7_R0_en),
    .W0_addr(mem_14_7_W0_addr),
    .W0_clk(mem_14_7_W0_clk),
    .W0_data(mem_14_7_W0_data),
    .W0_en(mem_14_7_W0_en),
    .W0_mask(mem_14_7_W0_mask)
  );
  split_mem_0_ext mem_15_0 (
    .R0_addr(mem_15_0_R0_addr),
    .R0_clk(mem_15_0_R0_clk),
    .R0_data(mem_15_0_R0_data),
    .R0_en(mem_15_0_R0_en),
    .W0_addr(mem_15_0_W0_addr),
    .W0_clk(mem_15_0_W0_clk),
    .W0_data(mem_15_0_W0_data),
    .W0_en(mem_15_0_W0_en),
    .W0_mask(mem_15_0_W0_mask)
  );
  split_mem_0_ext mem_15_1 (
    .R0_addr(mem_15_1_R0_addr),
    .R0_clk(mem_15_1_R0_clk),
    .R0_data(mem_15_1_R0_data),
    .R0_en(mem_15_1_R0_en),
    .W0_addr(mem_15_1_W0_addr),
    .W0_clk(mem_15_1_W0_clk),
    .W0_data(mem_15_1_W0_data),
    .W0_en(mem_15_1_W0_en),
    .W0_mask(mem_15_1_W0_mask)
  );
  split_mem_0_ext mem_15_2 (
    .R0_addr(mem_15_2_R0_addr),
    .R0_clk(mem_15_2_R0_clk),
    .R0_data(mem_15_2_R0_data),
    .R0_en(mem_15_2_R0_en),
    .W0_addr(mem_15_2_W0_addr),
    .W0_clk(mem_15_2_W0_clk),
    .W0_data(mem_15_2_W0_data),
    .W0_en(mem_15_2_W0_en),
    .W0_mask(mem_15_2_W0_mask)
  );
  split_mem_0_ext mem_15_3 (
    .R0_addr(mem_15_3_R0_addr),
    .R0_clk(mem_15_3_R0_clk),
    .R0_data(mem_15_3_R0_data),
    .R0_en(mem_15_3_R0_en),
    .W0_addr(mem_15_3_W0_addr),
    .W0_clk(mem_15_3_W0_clk),
    .W0_data(mem_15_3_W0_data),
    .W0_en(mem_15_3_W0_en),
    .W0_mask(mem_15_3_W0_mask)
  );
  split_mem_0_ext mem_15_4 (
    .R0_addr(mem_15_4_R0_addr),
    .R0_clk(mem_15_4_R0_clk),
    .R0_data(mem_15_4_R0_data),
    .R0_en(mem_15_4_R0_en),
    .W0_addr(mem_15_4_W0_addr),
    .W0_clk(mem_15_4_W0_clk),
    .W0_data(mem_15_4_W0_data),
    .W0_en(mem_15_4_W0_en),
    .W0_mask(mem_15_4_W0_mask)
  );
  split_mem_0_ext mem_15_5 (
    .R0_addr(mem_15_5_R0_addr),
    .R0_clk(mem_15_5_R0_clk),
    .R0_data(mem_15_5_R0_data),
    .R0_en(mem_15_5_R0_en),
    .W0_addr(mem_15_5_W0_addr),
    .W0_clk(mem_15_5_W0_clk),
    .W0_data(mem_15_5_W0_data),
    .W0_en(mem_15_5_W0_en),
    .W0_mask(mem_15_5_W0_mask)
  );
  split_mem_0_ext mem_15_6 (
    .R0_addr(mem_15_6_R0_addr),
    .R0_clk(mem_15_6_R0_clk),
    .R0_data(mem_15_6_R0_data),
    .R0_en(mem_15_6_R0_en),
    .W0_addr(mem_15_6_W0_addr),
    .W0_clk(mem_15_6_W0_clk),
    .W0_data(mem_15_6_W0_data),
    .W0_en(mem_15_6_W0_en),
    .W0_mask(mem_15_6_W0_mask)
  );
  split_mem_0_ext mem_15_7 (
    .R0_addr(mem_15_7_R0_addr),
    .R0_clk(mem_15_7_R0_clk),
    .R0_data(mem_15_7_R0_data),
    .R0_en(mem_15_7_R0_en),
    .W0_addr(mem_15_7_W0_addr),
    .W0_clk(mem_15_7_W0_clk),
    .W0_data(mem_15_7_W0_data),
    .W0_en(mem_15_7_W0_en),
    .W0_mask(mem_15_7_W0_mask)
  );
  split_mem_0_ext mem_16_0 (
    .R0_addr(mem_16_0_R0_addr),
    .R0_clk(mem_16_0_R0_clk),
    .R0_data(mem_16_0_R0_data),
    .R0_en(mem_16_0_R0_en),
    .W0_addr(mem_16_0_W0_addr),
    .W0_clk(mem_16_0_W0_clk),
    .W0_data(mem_16_0_W0_data),
    .W0_en(mem_16_0_W0_en),
    .W0_mask(mem_16_0_W0_mask)
  );
  split_mem_0_ext mem_16_1 (
    .R0_addr(mem_16_1_R0_addr),
    .R0_clk(mem_16_1_R0_clk),
    .R0_data(mem_16_1_R0_data),
    .R0_en(mem_16_1_R0_en),
    .W0_addr(mem_16_1_W0_addr),
    .W0_clk(mem_16_1_W0_clk),
    .W0_data(mem_16_1_W0_data),
    .W0_en(mem_16_1_W0_en),
    .W0_mask(mem_16_1_W0_mask)
  );
  split_mem_0_ext mem_16_2 (
    .R0_addr(mem_16_2_R0_addr),
    .R0_clk(mem_16_2_R0_clk),
    .R0_data(mem_16_2_R0_data),
    .R0_en(mem_16_2_R0_en),
    .W0_addr(mem_16_2_W0_addr),
    .W0_clk(mem_16_2_W0_clk),
    .W0_data(mem_16_2_W0_data),
    .W0_en(mem_16_2_W0_en),
    .W0_mask(mem_16_2_W0_mask)
  );
  split_mem_0_ext mem_16_3 (
    .R0_addr(mem_16_3_R0_addr),
    .R0_clk(mem_16_3_R0_clk),
    .R0_data(mem_16_3_R0_data),
    .R0_en(mem_16_3_R0_en),
    .W0_addr(mem_16_3_W0_addr),
    .W0_clk(mem_16_3_W0_clk),
    .W0_data(mem_16_3_W0_data),
    .W0_en(mem_16_3_W0_en),
    .W0_mask(mem_16_3_W0_mask)
  );
  split_mem_0_ext mem_16_4 (
    .R0_addr(mem_16_4_R0_addr),
    .R0_clk(mem_16_4_R0_clk),
    .R0_data(mem_16_4_R0_data),
    .R0_en(mem_16_4_R0_en),
    .W0_addr(mem_16_4_W0_addr),
    .W0_clk(mem_16_4_W0_clk),
    .W0_data(mem_16_4_W0_data),
    .W0_en(mem_16_4_W0_en),
    .W0_mask(mem_16_4_W0_mask)
  );
  split_mem_0_ext mem_16_5 (
    .R0_addr(mem_16_5_R0_addr),
    .R0_clk(mem_16_5_R0_clk),
    .R0_data(mem_16_5_R0_data),
    .R0_en(mem_16_5_R0_en),
    .W0_addr(mem_16_5_W0_addr),
    .W0_clk(mem_16_5_W0_clk),
    .W0_data(mem_16_5_W0_data),
    .W0_en(mem_16_5_W0_en),
    .W0_mask(mem_16_5_W0_mask)
  );
  split_mem_0_ext mem_16_6 (
    .R0_addr(mem_16_6_R0_addr),
    .R0_clk(mem_16_6_R0_clk),
    .R0_data(mem_16_6_R0_data),
    .R0_en(mem_16_6_R0_en),
    .W0_addr(mem_16_6_W0_addr),
    .W0_clk(mem_16_6_W0_clk),
    .W0_data(mem_16_6_W0_data),
    .W0_en(mem_16_6_W0_en),
    .W0_mask(mem_16_6_W0_mask)
  );
  split_mem_0_ext mem_16_7 (
    .R0_addr(mem_16_7_R0_addr),
    .R0_clk(mem_16_7_R0_clk),
    .R0_data(mem_16_7_R0_data),
    .R0_en(mem_16_7_R0_en),
    .W0_addr(mem_16_7_W0_addr),
    .W0_clk(mem_16_7_W0_clk),
    .W0_data(mem_16_7_W0_data),
    .W0_en(mem_16_7_W0_en),
    .W0_mask(mem_16_7_W0_mask)
  );
  split_mem_0_ext mem_17_0 (
    .R0_addr(mem_17_0_R0_addr),
    .R0_clk(mem_17_0_R0_clk),
    .R0_data(mem_17_0_R0_data),
    .R0_en(mem_17_0_R0_en),
    .W0_addr(mem_17_0_W0_addr),
    .W0_clk(mem_17_0_W0_clk),
    .W0_data(mem_17_0_W0_data),
    .W0_en(mem_17_0_W0_en),
    .W0_mask(mem_17_0_W0_mask)
  );
  split_mem_0_ext mem_17_1 (
    .R0_addr(mem_17_1_R0_addr),
    .R0_clk(mem_17_1_R0_clk),
    .R0_data(mem_17_1_R0_data),
    .R0_en(mem_17_1_R0_en),
    .W0_addr(mem_17_1_W0_addr),
    .W0_clk(mem_17_1_W0_clk),
    .W0_data(mem_17_1_W0_data),
    .W0_en(mem_17_1_W0_en),
    .W0_mask(mem_17_1_W0_mask)
  );
  split_mem_0_ext mem_17_2 (
    .R0_addr(mem_17_2_R0_addr),
    .R0_clk(mem_17_2_R0_clk),
    .R0_data(mem_17_2_R0_data),
    .R0_en(mem_17_2_R0_en),
    .W0_addr(mem_17_2_W0_addr),
    .W0_clk(mem_17_2_W0_clk),
    .W0_data(mem_17_2_W0_data),
    .W0_en(mem_17_2_W0_en),
    .W0_mask(mem_17_2_W0_mask)
  );
  split_mem_0_ext mem_17_3 (
    .R0_addr(mem_17_3_R0_addr),
    .R0_clk(mem_17_3_R0_clk),
    .R0_data(mem_17_3_R0_data),
    .R0_en(mem_17_3_R0_en),
    .W0_addr(mem_17_3_W0_addr),
    .W0_clk(mem_17_3_W0_clk),
    .W0_data(mem_17_3_W0_data),
    .W0_en(mem_17_3_W0_en),
    .W0_mask(mem_17_3_W0_mask)
  );
  split_mem_0_ext mem_17_4 (
    .R0_addr(mem_17_4_R0_addr),
    .R0_clk(mem_17_4_R0_clk),
    .R0_data(mem_17_4_R0_data),
    .R0_en(mem_17_4_R0_en),
    .W0_addr(mem_17_4_W0_addr),
    .W0_clk(mem_17_4_W0_clk),
    .W0_data(mem_17_4_W0_data),
    .W0_en(mem_17_4_W0_en),
    .W0_mask(mem_17_4_W0_mask)
  );
  split_mem_0_ext mem_17_5 (
    .R0_addr(mem_17_5_R0_addr),
    .R0_clk(mem_17_5_R0_clk),
    .R0_data(mem_17_5_R0_data),
    .R0_en(mem_17_5_R0_en),
    .W0_addr(mem_17_5_W0_addr),
    .W0_clk(mem_17_5_W0_clk),
    .W0_data(mem_17_5_W0_data),
    .W0_en(mem_17_5_W0_en),
    .W0_mask(mem_17_5_W0_mask)
  );
  split_mem_0_ext mem_17_6 (
    .R0_addr(mem_17_6_R0_addr),
    .R0_clk(mem_17_6_R0_clk),
    .R0_data(mem_17_6_R0_data),
    .R0_en(mem_17_6_R0_en),
    .W0_addr(mem_17_6_W0_addr),
    .W0_clk(mem_17_6_W0_clk),
    .W0_data(mem_17_6_W0_data),
    .W0_en(mem_17_6_W0_en),
    .W0_mask(mem_17_6_W0_mask)
  );
  split_mem_0_ext mem_17_7 (
    .R0_addr(mem_17_7_R0_addr),
    .R0_clk(mem_17_7_R0_clk),
    .R0_data(mem_17_7_R0_data),
    .R0_en(mem_17_7_R0_en),
    .W0_addr(mem_17_7_W0_addr),
    .W0_clk(mem_17_7_W0_clk),
    .W0_data(mem_17_7_W0_data),
    .W0_en(mem_17_7_W0_en),
    .W0_mask(mem_17_7_W0_mask)
  );
  split_mem_0_ext mem_18_0 (
    .R0_addr(mem_18_0_R0_addr),
    .R0_clk(mem_18_0_R0_clk),
    .R0_data(mem_18_0_R0_data),
    .R0_en(mem_18_0_R0_en),
    .W0_addr(mem_18_0_W0_addr),
    .W0_clk(mem_18_0_W0_clk),
    .W0_data(mem_18_0_W0_data),
    .W0_en(mem_18_0_W0_en),
    .W0_mask(mem_18_0_W0_mask)
  );
  split_mem_0_ext mem_18_1 (
    .R0_addr(mem_18_1_R0_addr),
    .R0_clk(mem_18_1_R0_clk),
    .R0_data(mem_18_1_R0_data),
    .R0_en(mem_18_1_R0_en),
    .W0_addr(mem_18_1_W0_addr),
    .W0_clk(mem_18_1_W0_clk),
    .W0_data(mem_18_1_W0_data),
    .W0_en(mem_18_1_W0_en),
    .W0_mask(mem_18_1_W0_mask)
  );
  split_mem_0_ext mem_18_2 (
    .R0_addr(mem_18_2_R0_addr),
    .R0_clk(mem_18_2_R0_clk),
    .R0_data(mem_18_2_R0_data),
    .R0_en(mem_18_2_R0_en),
    .W0_addr(mem_18_2_W0_addr),
    .W0_clk(mem_18_2_W0_clk),
    .W0_data(mem_18_2_W0_data),
    .W0_en(mem_18_2_W0_en),
    .W0_mask(mem_18_2_W0_mask)
  );
  split_mem_0_ext mem_18_3 (
    .R0_addr(mem_18_3_R0_addr),
    .R0_clk(mem_18_3_R0_clk),
    .R0_data(mem_18_3_R0_data),
    .R0_en(mem_18_3_R0_en),
    .W0_addr(mem_18_3_W0_addr),
    .W0_clk(mem_18_3_W0_clk),
    .W0_data(mem_18_3_W0_data),
    .W0_en(mem_18_3_W0_en),
    .W0_mask(mem_18_3_W0_mask)
  );
  split_mem_0_ext mem_18_4 (
    .R0_addr(mem_18_4_R0_addr),
    .R0_clk(mem_18_4_R0_clk),
    .R0_data(mem_18_4_R0_data),
    .R0_en(mem_18_4_R0_en),
    .W0_addr(mem_18_4_W0_addr),
    .W0_clk(mem_18_4_W0_clk),
    .W0_data(mem_18_4_W0_data),
    .W0_en(mem_18_4_W0_en),
    .W0_mask(mem_18_4_W0_mask)
  );
  split_mem_0_ext mem_18_5 (
    .R0_addr(mem_18_5_R0_addr),
    .R0_clk(mem_18_5_R0_clk),
    .R0_data(mem_18_5_R0_data),
    .R0_en(mem_18_5_R0_en),
    .W0_addr(mem_18_5_W0_addr),
    .W0_clk(mem_18_5_W0_clk),
    .W0_data(mem_18_5_W0_data),
    .W0_en(mem_18_5_W0_en),
    .W0_mask(mem_18_5_W0_mask)
  );
  split_mem_0_ext mem_18_6 (
    .R0_addr(mem_18_6_R0_addr),
    .R0_clk(mem_18_6_R0_clk),
    .R0_data(mem_18_6_R0_data),
    .R0_en(mem_18_6_R0_en),
    .W0_addr(mem_18_6_W0_addr),
    .W0_clk(mem_18_6_W0_clk),
    .W0_data(mem_18_6_W0_data),
    .W0_en(mem_18_6_W0_en),
    .W0_mask(mem_18_6_W0_mask)
  );
  split_mem_0_ext mem_18_7 (
    .R0_addr(mem_18_7_R0_addr),
    .R0_clk(mem_18_7_R0_clk),
    .R0_data(mem_18_7_R0_data),
    .R0_en(mem_18_7_R0_en),
    .W0_addr(mem_18_7_W0_addr),
    .W0_clk(mem_18_7_W0_clk),
    .W0_data(mem_18_7_W0_data),
    .W0_en(mem_18_7_W0_en),
    .W0_mask(mem_18_7_W0_mask)
  );
  split_mem_0_ext mem_19_0 (
    .R0_addr(mem_19_0_R0_addr),
    .R0_clk(mem_19_0_R0_clk),
    .R0_data(mem_19_0_R0_data),
    .R0_en(mem_19_0_R0_en),
    .W0_addr(mem_19_0_W0_addr),
    .W0_clk(mem_19_0_W0_clk),
    .W0_data(mem_19_0_W0_data),
    .W0_en(mem_19_0_W0_en),
    .W0_mask(mem_19_0_W0_mask)
  );
  split_mem_0_ext mem_19_1 (
    .R0_addr(mem_19_1_R0_addr),
    .R0_clk(mem_19_1_R0_clk),
    .R0_data(mem_19_1_R0_data),
    .R0_en(mem_19_1_R0_en),
    .W0_addr(mem_19_1_W0_addr),
    .W0_clk(mem_19_1_W0_clk),
    .W0_data(mem_19_1_W0_data),
    .W0_en(mem_19_1_W0_en),
    .W0_mask(mem_19_1_W0_mask)
  );
  split_mem_0_ext mem_19_2 (
    .R0_addr(mem_19_2_R0_addr),
    .R0_clk(mem_19_2_R0_clk),
    .R0_data(mem_19_2_R0_data),
    .R0_en(mem_19_2_R0_en),
    .W0_addr(mem_19_2_W0_addr),
    .W0_clk(mem_19_2_W0_clk),
    .W0_data(mem_19_2_W0_data),
    .W0_en(mem_19_2_W0_en),
    .W0_mask(mem_19_2_W0_mask)
  );
  split_mem_0_ext mem_19_3 (
    .R0_addr(mem_19_3_R0_addr),
    .R0_clk(mem_19_3_R0_clk),
    .R0_data(mem_19_3_R0_data),
    .R0_en(mem_19_3_R0_en),
    .W0_addr(mem_19_3_W0_addr),
    .W0_clk(mem_19_3_W0_clk),
    .W0_data(mem_19_3_W0_data),
    .W0_en(mem_19_3_W0_en),
    .W0_mask(mem_19_3_W0_mask)
  );
  split_mem_0_ext mem_19_4 (
    .R0_addr(mem_19_4_R0_addr),
    .R0_clk(mem_19_4_R0_clk),
    .R0_data(mem_19_4_R0_data),
    .R0_en(mem_19_4_R0_en),
    .W0_addr(mem_19_4_W0_addr),
    .W0_clk(mem_19_4_W0_clk),
    .W0_data(mem_19_4_W0_data),
    .W0_en(mem_19_4_W0_en),
    .W0_mask(mem_19_4_W0_mask)
  );
  split_mem_0_ext mem_19_5 (
    .R0_addr(mem_19_5_R0_addr),
    .R0_clk(mem_19_5_R0_clk),
    .R0_data(mem_19_5_R0_data),
    .R0_en(mem_19_5_R0_en),
    .W0_addr(mem_19_5_W0_addr),
    .W0_clk(mem_19_5_W0_clk),
    .W0_data(mem_19_5_W0_data),
    .W0_en(mem_19_5_W0_en),
    .W0_mask(mem_19_5_W0_mask)
  );
  split_mem_0_ext mem_19_6 (
    .R0_addr(mem_19_6_R0_addr),
    .R0_clk(mem_19_6_R0_clk),
    .R0_data(mem_19_6_R0_data),
    .R0_en(mem_19_6_R0_en),
    .W0_addr(mem_19_6_W0_addr),
    .W0_clk(mem_19_6_W0_clk),
    .W0_data(mem_19_6_W0_data),
    .W0_en(mem_19_6_W0_en),
    .W0_mask(mem_19_6_W0_mask)
  );
  split_mem_0_ext mem_19_7 (
    .R0_addr(mem_19_7_R0_addr),
    .R0_clk(mem_19_7_R0_clk),
    .R0_data(mem_19_7_R0_data),
    .R0_en(mem_19_7_R0_en),
    .W0_addr(mem_19_7_W0_addr),
    .W0_clk(mem_19_7_W0_clk),
    .W0_data(mem_19_7_W0_data),
    .W0_en(mem_19_7_W0_en),
    .W0_mask(mem_19_7_W0_mask)
  );
  split_mem_0_ext mem_20_0 (
    .R0_addr(mem_20_0_R0_addr),
    .R0_clk(mem_20_0_R0_clk),
    .R0_data(mem_20_0_R0_data),
    .R0_en(mem_20_0_R0_en),
    .W0_addr(mem_20_0_W0_addr),
    .W0_clk(mem_20_0_W0_clk),
    .W0_data(mem_20_0_W0_data),
    .W0_en(mem_20_0_W0_en),
    .W0_mask(mem_20_0_W0_mask)
  );
  split_mem_0_ext mem_20_1 (
    .R0_addr(mem_20_1_R0_addr),
    .R0_clk(mem_20_1_R0_clk),
    .R0_data(mem_20_1_R0_data),
    .R0_en(mem_20_1_R0_en),
    .W0_addr(mem_20_1_W0_addr),
    .W0_clk(mem_20_1_W0_clk),
    .W0_data(mem_20_1_W0_data),
    .W0_en(mem_20_1_W0_en),
    .W0_mask(mem_20_1_W0_mask)
  );
  split_mem_0_ext mem_20_2 (
    .R0_addr(mem_20_2_R0_addr),
    .R0_clk(mem_20_2_R0_clk),
    .R0_data(mem_20_2_R0_data),
    .R0_en(mem_20_2_R0_en),
    .W0_addr(mem_20_2_W0_addr),
    .W0_clk(mem_20_2_W0_clk),
    .W0_data(mem_20_2_W0_data),
    .W0_en(mem_20_2_W0_en),
    .W0_mask(mem_20_2_W0_mask)
  );
  split_mem_0_ext mem_20_3 (
    .R0_addr(mem_20_3_R0_addr),
    .R0_clk(mem_20_3_R0_clk),
    .R0_data(mem_20_3_R0_data),
    .R0_en(mem_20_3_R0_en),
    .W0_addr(mem_20_3_W0_addr),
    .W0_clk(mem_20_3_W0_clk),
    .W0_data(mem_20_3_W0_data),
    .W0_en(mem_20_3_W0_en),
    .W0_mask(mem_20_3_W0_mask)
  );
  split_mem_0_ext mem_20_4 (
    .R0_addr(mem_20_4_R0_addr),
    .R0_clk(mem_20_4_R0_clk),
    .R0_data(mem_20_4_R0_data),
    .R0_en(mem_20_4_R0_en),
    .W0_addr(mem_20_4_W0_addr),
    .W0_clk(mem_20_4_W0_clk),
    .W0_data(mem_20_4_W0_data),
    .W0_en(mem_20_4_W0_en),
    .W0_mask(mem_20_4_W0_mask)
  );
  split_mem_0_ext mem_20_5 (
    .R0_addr(mem_20_5_R0_addr),
    .R0_clk(mem_20_5_R0_clk),
    .R0_data(mem_20_5_R0_data),
    .R0_en(mem_20_5_R0_en),
    .W0_addr(mem_20_5_W0_addr),
    .W0_clk(mem_20_5_W0_clk),
    .W0_data(mem_20_5_W0_data),
    .W0_en(mem_20_5_W0_en),
    .W0_mask(mem_20_5_W0_mask)
  );
  split_mem_0_ext mem_20_6 (
    .R0_addr(mem_20_6_R0_addr),
    .R0_clk(mem_20_6_R0_clk),
    .R0_data(mem_20_6_R0_data),
    .R0_en(mem_20_6_R0_en),
    .W0_addr(mem_20_6_W0_addr),
    .W0_clk(mem_20_6_W0_clk),
    .W0_data(mem_20_6_W0_data),
    .W0_en(mem_20_6_W0_en),
    .W0_mask(mem_20_6_W0_mask)
  );
  split_mem_0_ext mem_20_7 (
    .R0_addr(mem_20_7_R0_addr),
    .R0_clk(mem_20_7_R0_clk),
    .R0_data(mem_20_7_R0_data),
    .R0_en(mem_20_7_R0_en),
    .W0_addr(mem_20_7_W0_addr),
    .W0_clk(mem_20_7_W0_clk),
    .W0_data(mem_20_7_W0_data),
    .W0_en(mem_20_7_W0_en),
    .W0_mask(mem_20_7_W0_mask)
  );
  split_mem_0_ext mem_21_0 (
    .R0_addr(mem_21_0_R0_addr),
    .R0_clk(mem_21_0_R0_clk),
    .R0_data(mem_21_0_R0_data),
    .R0_en(mem_21_0_R0_en),
    .W0_addr(mem_21_0_W0_addr),
    .W0_clk(mem_21_0_W0_clk),
    .W0_data(mem_21_0_W0_data),
    .W0_en(mem_21_0_W0_en),
    .W0_mask(mem_21_0_W0_mask)
  );
  split_mem_0_ext mem_21_1 (
    .R0_addr(mem_21_1_R0_addr),
    .R0_clk(mem_21_1_R0_clk),
    .R0_data(mem_21_1_R0_data),
    .R0_en(mem_21_1_R0_en),
    .W0_addr(mem_21_1_W0_addr),
    .W0_clk(mem_21_1_W0_clk),
    .W0_data(mem_21_1_W0_data),
    .W0_en(mem_21_1_W0_en),
    .W0_mask(mem_21_1_W0_mask)
  );
  split_mem_0_ext mem_21_2 (
    .R0_addr(mem_21_2_R0_addr),
    .R0_clk(mem_21_2_R0_clk),
    .R0_data(mem_21_2_R0_data),
    .R0_en(mem_21_2_R0_en),
    .W0_addr(mem_21_2_W0_addr),
    .W0_clk(mem_21_2_W0_clk),
    .W0_data(mem_21_2_W0_data),
    .W0_en(mem_21_2_W0_en),
    .W0_mask(mem_21_2_W0_mask)
  );
  split_mem_0_ext mem_21_3 (
    .R0_addr(mem_21_3_R0_addr),
    .R0_clk(mem_21_3_R0_clk),
    .R0_data(mem_21_3_R0_data),
    .R0_en(mem_21_3_R0_en),
    .W0_addr(mem_21_3_W0_addr),
    .W0_clk(mem_21_3_W0_clk),
    .W0_data(mem_21_3_W0_data),
    .W0_en(mem_21_3_W0_en),
    .W0_mask(mem_21_3_W0_mask)
  );
  split_mem_0_ext mem_21_4 (
    .R0_addr(mem_21_4_R0_addr),
    .R0_clk(mem_21_4_R0_clk),
    .R0_data(mem_21_4_R0_data),
    .R0_en(mem_21_4_R0_en),
    .W0_addr(mem_21_4_W0_addr),
    .W0_clk(mem_21_4_W0_clk),
    .W0_data(mem_21_4_W0_data),
    .W0_en(mem_21_4_W0_en),
    .W0_mask(mem_21_4_W0_mask)
  );
  split_mem_0_ext mem_21_5 (
    .R0_addr(mem_21_5_R0_addr),
    .R0_clk(mem_21_5_R0_clk),
    .R0_data(mem_21_5_R0_data),
    .R0_en(mem_21_5_R0_en),
    .W0_addr(mem_21_5_W0_addr),
    .W0_clk(mem_21_5_W0_clk),
    .W0_data(mem_21_5_W0_data),
    .W0_en(mem_21_5_W0_en),
    .W0_mask(mem_21_5_W0_mask)
  );
  split_mem_0_ext mem_21_6 (
    .R0_addr(mem_21_6_R0_addr),
    .R0_clk(mem_21_6_R0_clk),
    .R0_data(mem_21_6_R0_data),
    .R0_en(mem_21_6_R0_en),
    .W0_addr(mem_21_6_W0_addr),
    .W0_clk(mem_21_6_W0_clk),
    .W0_data(mem_21_6_W0_data),
    .W0_en(mem_21_6_W0_en),
    .W0_mask(mem_21_6_W0_mask)
  );
  split_mem_0_ext mem_21_7 (
    .R0_addr(mem_21_7_R0_addr),
    .R0_clk(mem_21_7_R0_clk),
    .R0_data(mem_21_7_R0_data),
    .R0_en(mem_21_7_R0_en),
    .W0_addr(mem_21_7_W0_addr),
    .W0_clk(mem_21_7_W0_clk),
    .W0_data(mem_21_7_W0_data),
    .W0_en(mem_21_7_W0_en),
    .W0_mask(mem_21_7_W0_mask)
  );
  split_mem_0_ext mem_22_0 (
    .R0_addr(mem_22_0_R0_addr),
    .R0_clk(mem_22_0_R0_clk),
    .R0_data(mem_22_0_R0_data),
    .R0_en(mem_22_0_R0_en),
    .W0_addr(mem_22_0_W0_addr),
    .W0_clk(mem_22_0_W0_clk),
    .W0_data(mem_22_0_W0_data),
    .W0_en(mem_22_0_W0_en),
    .W0_mask(mem_22_0_W0_mask)
  );
  split_mem_0_ext mem_22_1 (
    .R0_addr(mem_22_1_R0_addr),
    .R0_clk(mem_22_1_R0_clk),
    .R0_data(mem_22_1_R0_data),
    .R0_en(mem_22_1_R0_en),
    .W0_addr(mem_22_1_W0_addr),
    .W0_clk(mem_22_1_W0_clk),
    .W0_data(mem_22_1_W0_data),
    .W0_en(mem_22_1_W0_en),
    .W0_mask(mem_22_1_W0_mask)
  );
  split_mem_0_ext mem_22_2 (
    .R0_addr(mem_22_2_R0_addr),
    .R0_clk(mem_22_2_R0_clk),
    .R0_data(mem_22_2_R0_data),
    .R0_en(mem_22_2_R0_en),
    .W0_addr(mem_22_2_W0_addr),
    .W0_clk(mem_22_2_W0_clk),
    .W0_data(mem_22_2_W0_data),
    .W0_en(mem_22_2_W0_en),
    .W0_mask(mem_22_2_W0_mask)
  );
  split_mem_0_ext mem_22_3 (
    .R0_addr(mem_22_3_R0_addr),
    .R0_clk(mem_22_3_R0_clk),
    .R0_data(mem_22_3_R0_data),
    .R0_en(mem_22_3_R0_en),
    .W0_addr(mem_22_3_W0_addr),
    .W0_clk(mem_22_3_W0_clk),
    .W0_data(mem_22_3_W0_data),
    .W0_en(mem_22_3_W0_en),
    .W0_mask(mem_22_3_W0_mask)
  );
  split_mem_0_ext mem_22_4 (
    .R0_addr(mem_22_4_R0_addr),
    .R0_clk(mem_22_4_R0_clk),
    .R0_data(mem_22_4_R0_data),
    .R0_en(mem_22_4_R0_en),
    .W0_addr(mem_22_4_W0_addr),
    .W0_clk(mem_22_4_W0_clk),
    .W0_data(mem_22_4_W0_data),
    .W0_en(mem_22_4_W0_en),
    .W0_mask(mem_22_4_W0_mask)
  );
  split_mem_0_ext mem_22_5 (
    .R0_addr(mem_22_5_R0_addr),
    .R0_clk(mem_22_5_R0_clk),
    .R0_data(mem_22_5_R0_data),
    .R0_en(mem_22_5_R0_en),
    .W0_addr(mem_22_5_W0_addr),
    .W0_clk(mem_22_5_W0_clk),
    .W0_data(mem_22_5_W0_data),
    .W0_en(mem_22_5_W0_en),
    .W0_mask(mem_22_5_W0_mask)
  );
  split_mem_0_ext mem_22_6 (
    .R0_addr(mem_22_6_R0_addr),
    .R0_clk(mem_22_6_R0_clk),
    .R0_data(mem_22_6_R0_data),
    .R0_en(mem_22_6_R0_en),
    .W0_addr(mem_22_6_W0_addr),
    .W0_clk(mem_22_6_W0_clk),
    .W0_data(mem_22_6_W0_data),
    .W0_en(mem_22_6_W0_en),
    .W0_mask(mem_22_6_W0_mask)
  );
  split_mem_0_ext mem_22_7 (
    .R0_addr(mem_22_7_R0_addr),
    .R0_clk(mem_22_7_R0_clk),
    .R0_data(mem_22_7_R0_data),
    .R0_en(mem_22_7_R0_en),
    .W0_addr(mem_22_7_W0_addr),
    .W0_clk(mem_22_7_W0_clk),
    .W0_data(mem_22_7_W0_data),
    .W0_en(mem_22_7_W0_en),
    .W0_mask(mem_22_7_W0_mask)
  );
  split_mem_0_ext mem_23_0 (
    .R0_addr(mem_23_0_R0_addr),
    .R0_clk(mem_23_0_R0_clk),
    .R0_data(mem_23_0_R0_data),
    .R0_en(mem_23_0_R0_en),
    .W0_addr(mem_23_0_W0_addr),
    .W0_clk(mem_23_0_W0_clk),
    .W0_data(mem_23_0_W0_data),
    .W0_en(mem_23_0_W0_en),
    .W0_mask(mem_23_0_W0_mask)
  );
  split_mem_0_ext mem_23_1 (
    .R0_addr(mem_23_1_R0_addr),
    .R0_clk(mem_23_1_R0_clk),
    .R0_data(mem_23_1_R0_data),
    .R0_en(mem_23_1_R0_en),
    .W0_addr(mem_23_1_W0_addr),
    .W0_clk(mem_23_1_W0_clk),
    .W0_data(mem_23_1_W0_data),
    .W0_en(mem_23_1_W0_en),
    .W0_mask(mem_23_1_W0_mask)
  );
  split_mem_0_ext mem_23_2 (
    .R0_addr(mem_23_2_R0_addr),
    .R0_clk(mem_23_2_R0_clk),
    .R0_data(mem_23_2_R0_data),
    .R0_en(mem_23_2_R0_en),
    .W0_addr(mem_23_2_W0_addr),
    .W0_clk(mem_23_2_W0_clk),
    .W0_data(mem_23_2_W0_data),
    .W0_en(mem_23_2_W0_en),
    .W0_mask(mem_23_2_W0_mask)
  );
  split_mem_0_ext mem_23_3 (
    .R0_addr(mem_23_3_R0_addr),
    .R0_clk(mem_23_3_R0_clk),
    .R0_data(mem_23_3_R0_data),
    .R0_en(mem_23_3_R0_en),
    .W0_addr(mem_23_3_W0_addr),
    .W0_clk(mem_23_3_W0_clk),
    .W0_data(mem_23_3_W0_data),
    .W0_en(mem_23_3_W0_en),
    .W0_mask(mem_23_3_W0_mask)
  );
  split_mem_0_ext mem_23_4 (
    .R0_addr(mem_23_4_R0_addr),
    .R0_clk(mem_23_4_R0_clk),
    .R0_data(mem_23_4_R0_data),
    .R0_en(mem_23_4_R0_en),
    .W0_addr(mem_23_4_W0_addr),
    .W0_clk(mem_23_4_W0_clk),
    .W0_data(mem_23_4_W0_data),
    .W0_en(mem_23_4_W0_en),
    .W0_mask(mem_23_4_W0_mask)
  );
  split_mem_0_ext mem_23_5 (
    .R0_addr(mem_23_5_R0_addr),
    .R0_clk(mem_23_5_R0_clk),
    .R0_data(mem_23_5_R0_data),
    .R0_en(mem_23_5_R0_en),
    .W0_addr(mem_23_5_W0_addr),
    .W0_clk(mem_23_5_W0_clk),
    .W0_data(mem_23_5_W0_data),
    .W0_en(mem_23_5_W0_en),
    .W0_mask(mem_23_5_W0_mask)
  );
  split_mem_0_ext mem_23_6 (
    .R0_addr(mem_23_6_R0_addr),
    .R0_clk(mem_23_6_R0_clk),
    .R0_data(mem_23_6_R0_data),
    .R0_en(mem_23_6_R0_en),
    .W0_addr(mem_23_6_W0_addr),
    .W0_clk(mem_23_6_W0_clk),
    .W0_data(mem_23_6_W0_data),
    .W0_en(mem_23_6_W0_en),
    .W0_mask(mem_23_6_W0_mask)
  );
  split_mem_0_ext mem_23_7 (
    .R0_addr(mem_23_7_R0_addr),
    .R0_clk(mem_23_7_R0_clk),
    .R0_data(mem_23_7_R0_data),
    .R0_en(mem_23_7_R0_en),
    .W0_addr(mem_23_7_W0_addr),
    .W0_clk(mem_23_7_W0_clk),
    .W0_data(mem_23_7_W0_data),
    .W0_en(mem_23_7_W0_en),
    .W0_mask(mem_23_7_W0_mask)
  );
  split_mem_0_ext mem_24_0 (
    .R0_addr(mem_24_0_R0_addr),
    .R0_clk(mem_24_0_R0_clk),
    .R0_data(mem_24_0_R0_data),
    .R0_en(mem_24_0_R0_en),
    .W0_addr(mem_24_0_W0_addr),
    .W0_clk(mem_24_0_W0_clk),
    .W0_data(mem_24_0_W0_data),
    .W0_en(mem_24_0_W0_en),
    .W0_mask(mem_24_0_W0_mask)
  );
  split_mem_0_ext mem_24_1 (
    .R0_addr(mem_24_1_R0_addr),
    .R0_clk(mem_24_1_R0_clk),
    .R0_data(mem_24_1_R0_data),
    .R0_en(mem_24_1_R0_en),
    .W0_addr(mem_24_1_W0_addr),
    .W0_clk(mem_24_1_W0_clk),
    .W0_data(mem_24_1_W0_data),
    .W0_en(mem_24_1_W0_en),
    .W0_mask(mem_24_1_W0_mask)
  );
  split_mem_0_ext mem_24_2 (
    .R0_addr(mem_24_2_R0_addr),
    .R0_clk(mem_24_2_R0_clk),
    .R0_data(mem_24_2_R0_data),
    .R0_en(mem_24_2_R0_en),
    .W0_addr(mem_24_2_W0_addr),
    .W0_clk(mem_24_2_W0_clk),
    .W0_data(mem_24_2_W0_data),
    .W0_en(mem_24_2_W0_en),
    .W0_mask(mem_24_2_W0_mask)
  );
  split_mem_0_ext mem_24_3 (
    .R0_addr(mem_24_3_R0_addr),
    .R0_clk(mem_24_3_R0_clk),
    .R0_data(mem_24_3_R0_data),
    .R0_en(mem_24_3_R0_en),
    .W0_addr(mem_24_3_W0_addr),
    .W0_clk(mem_24_3_W0_clk),
    .W0_data(mem_24_3_W0_data),
    .W0_en(mem_24_3_W0_en),
    .W0_mask(mem_24_3_W0_mask)
  );
  split_mem_0_ext mem_24_4 (
    .R0_addr(mem_24_4_R0_addr),
    .R0_clk(mem_24_4_R0_clk),
    .R0_data(mem_24_4_R0_data),
    .R0_en(mem_24_4_R0_en),
    .W0_addr(mem_24_4_W0_addr),
    .W0_clk(mem_24_4_W0_clk),
    .W0_data(mem_24_4_W0_data),
    .W0_en(mem_24_4_W0_en),
    .W0_mask(mem_24_4_W0_mask)
  );
  split_mem_0_ext mem_24_5 (
    .R0_addr(mem_24_5_R0_addr),
    .R0_clk(mem_24_5_R0_clk),
    .R0_data(mem_24_5_R0_data),
    .R0_en(mem_24_5_R0_en),
    .W0_addr(mem_24_5_W0_addr),
    .W0_clk(mem_24_5_W0_clk),
    .W0_data(mem_24_5_W0_data),
    .W0_en(mem_24_5_W0_en),
    .W0_mask(mem_24_5_W0_mask)
  );
  split_mem_0_ext mem_24_6 (
    .R0_addr(mem_24_6_R0_addr),
    .R0_clk(mem_24_6_R0_clk),
    .R0_data(mem_24_6_R0_data),
    .R0_en(mem_24_6_R0_en),
    .W0_addr(mem_24_6_W0_addr),
    .W0_clk(mem_24_6_W0_clk),
    .W0_data(mem_24_6_W0_data),
    .W0_en(mem_24_6_W0_en),
    .W0_mask(mem_24_6_W0_mask)
  );
  split_mem_0_ext mem_24_7 (
    .R0_addr(mem_24_7_R0_addr),
    .R0_clk(mem_24_7_R0_clk),
    .R0_data(mem_24_7_R0_data),
    .R0_en(mem_24_7_R0_en),
    .W0_addr(mem_24_7_W0_addr),
    .W0_clk(mem_24_7_W0_clk),
    .W0_data(mem_24_7_W0_data),
    .W0_en(mem_24_7_W0_en),
    .W0_mask(mem_24_7_W0_mask)
  );
  split_mem_0_ext mem_25_0 (
    .R0_addr(mem_25_0_R0_addr),
    .R0_clk(mem_25_0_R0_clk),
    .R0_data(mem_25_0_R0_data),
    .R0_en(mem_25_0_R0_en),
    .W0_addr(mem_25_0_W0_addr),
    .W0_clk(mem_25_0_W0_clk),
    .W0_data(mem_25_0_W0_data),
    .W0_en(mem_25_0_W0_en),
    .W0_mask(mem_25_0_W0_mask)
  );
  split_mem_0_ext mem_25_1 (
    .R0_addr(mem_25_1_R0_addr),
    .R0_clk(mem_25_1_R0_clk),
    .R0_data(mem_25_1_R0_data),
    .R0_en(mem_25_1_R0_en),
    .W0_addr(mem_25_1_W0_addr),
    .W0_clk(mem_25_1_W0_clk),
    .W0_data(mem_25_1_W0_data),
    .W0_en(mem_25_1_W0_en),
    .W0_mask(mem_25_1_W0_mask)
  );
  split_mem_0_ext mem_25_2 (
    .R0_addr(mem_25_2_R0_addr),
    .R0_clk(mem_25_2_R0_clk),
    .R0_data(mem_25_2_R0_data),
    .R0_en(mem_25_2_R0_en),
    .W0_addr(mem_25_2_W0_addr),
    .W0_clk(mem_25_2_W0_clk),
    .W0_data(mem_25_2_W0_data),
    .W0_en(mem_25_2_W0_en),
    .W0_mask(mem_25_2_W0_mask)
  );
  split_mem_0_ext mem_25_3 (
    .R0_addr(mem_25_3_R0_addr),
    .R0_clk(mem_25_3_R0_clk),
    .R0_data(mem_25_3_R0_data),
    .R0_en(mem_25_3_R0_en),
    .W0_addr(mem_25_3_W0_addr),
    .W0_clk(mem_25_3_W0_clk),
    .W0_data(mem_25_3_W0_data),
    .W0_en(mem_25_3_W0_en),
    .W0_mask(mem_25_3_W0_mask)
  );
  split_mem_0_ext mem_25_4 (
    .R0_addr(mem_25_4_R0_addr),
    .R0_clk(mem_25_4_R0_clk),
    .R0_data(mem_25_4_R0_data),
    .R0_en(mem_25_4_R0_en),
    .W0_addr(mem_25_4_W0_addr),
    .W0_clk(mem_25_4_W0_clk),
    .W0_data(mem_25_4_W0_data),
    .W0_en(mem_25_4_W0_en),
    .W0_mask(mem_25_4_W0_mask)
  );
  split_mem_0_ext mem_25_5 (
    .R0_addr(mem_25_5_R0_addr),
    .R0_clk(mem_25_5_R0_clk),
    .R0_data(mem_25_5_R0_data),
    .R0_en(mem_25_5_R0_en),
    .W0_addr(mem_25_5_W0_addr),
    .W0_clk(mem_25_5_W0_clk),
    .W0_data(mem_25_5_W0_data),
    .W0_en(mem_25_5_W0_en),
    .W0_mask(mem_25_5_W0_mask)
  );
  split_mem_0_ext mem_25_6 (
    .R0_addr(mem_25_6_R0_addr),
    .R0_clk(mem_25_6_R0_clk),
    .R0_data(mem_25_6_R0_data),
    .R0_en(mem_25_6_R0_en),
    .W0_addr(mem_25_6_W0_addr),
    .W0_clk(mem_25_6_W0_clk),
    .W0_data(mem_25_6_W0_data),
    .W0_en(mem_25_6_W0_en),
    .W0_mask(mem_25_6_W0_mask)
  );
  split_mem_0_ext mem_25_7 (
    .R0_addr(mem_25_7_R0_addr),
    .R0_clk(mem_25_7_R0_clk),
    .R0_data(mem_25_7_R0_data),
    .R0_en(mem_25_7_R0_en),
    .W0_addr(mem_25_7_W0_addr),
    .W0_clk(mem_25_7_W0_clk),
    .W0_data(mem_25_7_W0_data),
    .W0_en(mem_25_7_W0_en),
    .W0_mask(mem_25_7_W0_mask)
  );
  split_mem_0_ext mem_26_0 (
    .R0_addr(mem_26_0_R0_addr),
    .R0_clk(mem_26_0_R0_clk),
    .R0_data(mem_26_0_R0_data),
    .R0_en(mem_26_0_R0_en),
    .W0_addr(mem_26_0_W0_addr),
    .W0_clk(mem_26_0_W0_clk),
    .W0_data(mem_26_0_W0_data),
    .W0_en(mem_26_0_W0_en),
    .W0_mask(mem_26_0_W0_mask)
  );
  split_mem_0_ext mem_26_1 (
    .R0_addr(mem_26_1_R0_addr),
    .R0_clk(mem_26_1_R0_clk),
    .R0_data(mem_26_1_R0_data),
    .R0_en(mem_26_1_R0_en),
    .W0_addr(mem_26_1_W0_addr),
    .W0_clk(mem_26_1_W0_clk),
    .W0_data(mem_26_1_W0_data),
    .W0_en(mem_26_1_W0_en),
    .W0_mask(mem_26_1_W0_mask)
  );
  split_mem_0_ext mem_26_2 (
    .R0_addr(mem_26_2_R0_addr),
    .R0_clk(mem_26_2_R0_clk),
    .R0_data(mem_26_2_R0_data),
    .R0_en(mem_26_2_R0_en),
    .W0_addr(mem_26_2_W0_addr),
    .W0_clk(mem_26_2_W0_clk),
    .W0_data(mem_26_2_W0_data),
    .W0_en(mem_26_2_W0_en),
    .W0_mask(mem_26_2_W0_mask)
  );
  split_mem_0_ext mem_26_3 (
    .R0_addr(mem_26_3_R0_addr),
    .R0_clk(mem_26_3_R0_clk),
    .R0_data(mem_26_3_R0_data),
    .R0_en(mem_26_3_R0_en),
    .W0_addr(mem_26_3_W0_addr),
    .W0_clk(mem_26_3_W0_clk),
    .W0_data(mem_26_3_W0_data),
    .W0_en(mem_26_3_W0_en),
    .W0_mask(mem_26_3_W0_mask)
  );
  split_mem_0_ext mem_26_4 (
    .R0_addr(mem_26_4_R0_addr),
    .R0_clk(mem_26_4_R0_clk),
    .R0_data(mem_26_4_R0_data),
    .R0_en(mem_26_4_R0_en),
    .W0_addr(mem_26_4_W0_addr),
    .W0_clk(mem_26_4_W0_clk),
    .W0_data(mem_26_4_W0_data),
    .W0_en(mem_26_4_W0_en),
    .W0_mask(mem_26_4_W0_mask)
  );
  split_mem_0_ext mem_26_5 (
    .R0_addr(mem_26_5_R0_addr),
    .R0_clk(mem_26_5_R0_clk),
    .R0_data(mem_26_5_R0_data),
    .R0_en(mem_26_5_R0_en),
    .W0_addr(mem_26_5_W0_addr),
    .W0_clk(mem_26_5_W0_clk),
    .W0_data(mem_26_5_W0_data),
    .W0_en(mem_26_5_W0_en),
    .W0_mask(mem_26_5_W0_mask)
  );
  split_mem_0_ext mem_26_6 (
    .R0_addr(mem_26_6_R0_addr),
    .R0_clk(mem_26_6_R0_clk),
    .R0_data(mem_26_6_R0_data),
    .R0_en(mem_26_6_R0_en),
    .W0_addr(mem_26_6_W0_addr),
    .W0_clk(mem_26_6_W0_clk),
    .W0_data(mem_26_6_W0_data),
    .W0_en(mem_26_6_W0_en),
    .W0_mask(mem_26_6_W0_mask)
  );
  split_mem_0_ext mem_26_7 (
    .R0_addr(mem_26_7_R0_addr),
    .R0_clk(mem_26_7_R0_clk),
    .R0_data(mem_26_7_R0_data),
    .R0_en(mem_26_7_R0_en),
    .W0_addr(mem_26_7_W0_addr),
    .W0_clk(mem_26_7_W0_clk),
    .W0_data(mem_26_7_W0_data),
    .W0_en(mem_26_7_W0_en),
    .W0_mask(mem_26_7_W0_mask)
  );
  split_mem_0_ext mem_27_0 (
    .R0_addr(mem_27_0_R0_addr),
    .R0_clk(mem_27_0_R0_clk),
    .R0_data(mem_27_0_R0_data),
    .R0_en(mem_27_0_R0_en),
    .W0_addr(mem_27_0_W0_addr),
    .W0_clk(mem_27_0_W0_clk),
    .W0_data(mem_27_0_W0_data),
    .W0_en(mem_27_0_W0_en),
    .W0_mask(mem_27_0_W0_mask)
  );
  split_mem_0_ext mem_27_1 (
    .R0_addr(mem_27_1_R0_addr),
    .R0_clk(mem_27_1_R0_clk),
    .R0_data(mem_27_1_R0_data),
    .R0_en(mem_27_1_R0_en),
    .W0_addr(mem_27_1_W0_addr),
    .W0_clk(mem_27_1_W0_clk),
    .W0_data(mem_27_1_W0_data),
    .W0_en(mem_27_1_W0_en),
    .W0_mask(mem_27_1_W0_mask)
  );
  split_mem_0_ext mem_27_2 (
    .R0_addr(mem_27_2_R0_addr),
    .R0_clk(mem_27_2_R0_clk),
    .R0_data(mem_27_2_R0_data),
    .R0_en(mem_27_2_R0_en),
    .W0_addr(mem_27_2_W0_addr),
    .W0_clk(mem_27_2_W0_clk),
    .W0_data(mem_27_2_W0_data),
    .W0_en(mem_27_2_W0_en),
    .W0_mask(mem_27_2_W0_mask)
  );
  split_mem_0_ext mem_27_3 (
    .R0_addr(mem_27_3_R0_addr),
    .R0_clk(mem_27_3_R0_clk),
    .R0_data(mem_27_3_R0_data),
    .R0_en(mem_27_3_R0_en),
    .W0_addr(mem_27_3_W0_addr),
    .W0_clk(mem_27_3_W0_clk),
    .W0_data(mem_27_3_W0_data),
    .W0_en(mem_27_3_W0_en),
    .W0_mask(mem_27_3_W0_mask)
  );
  split_mem_0_ext mem_27_4 (
    .R0_addr(mem_27_4_R0_addr),
    .R0_clk(mem_27_4_R0_clk),
    .R0_data(mem_27_4_R0_data),
    .R0_en(mem_27_4_R0_en),
    .W0_addr(mem_27_4_W0_addr),
    .W0_clk(mem_27_4_W0_clk),
    .W0_data(mem_27_4_W0_data),
    .W0_en(mem_27_4_W0_en),
    .W0_mask(mem_27_4_W0_mask)
  );
  split_mem_0_ext mem_27_5 (
    .R0_addr(mem_27_5_R0_addr),
    .R0_clk(mem_27_5_R0_clk),
    .R0_data(mem_27_5_R0_data),
    .R0_en(mem_27_5_R0_en),
    .W0_addr(mem_27_5_W0_addr),
    .W0_clk(mem_27_5_W0_clk),
    .W0_data(mem_27_5_W0_data),
    .W0_en(mem_27_5_W0_en),
    .W0_mask(mem_27_5_W0_mask)
  );
  split_mem_0_ext mem_27_6 (
    .R0_addr(mem_27_6_R0_addr),
    .R0_clk(mem_27_6_R0_clk),
    .R0_data(mem_27_6_R0_data),
    .R0_en(mem_27_6_R0_en),
    .W0_addr(mem_27_6_W0_addr),
    .W0_clk(mem_27_6_W0_clk),
    .W0_data(mem_27_6_W0_data),
    .W0_en(mem_27_6_W0_en),
    .W0_mask(mem_27_6_W0_mask)
  );
  split_mem_0_ext mem_27_7 (
    .R0_addr(mem_27_7_R0_addr),
    .R0_clk(mem_27_7_R0_clk),
    .R0_data(mem_27_7_R0_data),
    .R0_en(mem_27_7_R0_en),
    .W0_addr(mem_27_7_W0_addr),
    .W0_clk(mem_27_7_W0_clk),
    .W0_data(mem_27_7_W0_data),
    .W0_en(mem_27_7_W0_en),
    .W0_mask(mem_27_7_W0_mask)
  );
  split_mem_0_ext mem_28_0 (
    .R0_addr(mem_28_0_R0_addr),
    .R0_clk(mem_28_0_R0_clk),
    .R0_data(mem_28_0_R0_data),
    .R0_en(mem_28_0_R0_en),
    .W0_addr(mem_28_0_W0_addr),
    .W0_clk(mem_28_0_W0_clk),
    .W0_data(mem_28_0_W0_data),
    .W0_en(mem_28_0_W0_en),
    .W0_mask(mem_28_0_W0_mask)
  );
  split_mem_0_ext mem_28_1 (
    .R0_addr(mem_28_1_R0_addr),
    .R0_clk(mem_28_1_R0_clk),
    .R0_data(mem_28_1_R0_data),
    .R0_en(mem_28_1_R0_en),
    .W0_addr(mem_28_1_W0_addr),
    .W0_clk(mem_28_1_W0_clk),
    .W0_data(mem_28_1_W0_data),
    .W0_en(mem_28_1_W0_en),
    .W0_mask(mem_28_1_W0_mask)
  );
  split_mem_0_ext mem_28_2 (
    .R0_addr(mem_28_2_R0_addr),
    .R0_clk(mem_28_2_R0_clk),
    .R0_data(mem_28_2_R0_data),
    .R0_en(mem_28_2_R0_en),
    .W0_addr(mem_28_2_W0_addr),
    .W0_clk(mem_28_2_W0_clk),
    .W0_data(mem_28_2_W0_data),
    .W0_en(mem_28_2_W0_en),
    .W0_mask(mem_28_2_W0_mask)
  );
  split_mem_0_ext mem_28_3 (
    .R0_addr(mem_28_3_R0_addr),
    .R0_clk(mem_28_3_R0_clk),
    .R0_data(mem_28_3_R0_data),
    .R0_en(mem_28_3_R0_en),
    .W0_addr(mem_28_3_W0_addr),
    .W0_clk(mem_28_3_W0_clk),
    .W0_data(mem_28_3_W0_data),
    .W0_en(mem_28_3_W0_en),
    .W0_mask(mem_28_3_W0_mask)
  );
  split_mem_0_ext mem_28_4 (
    .R0_addr(mem_28_4_R0_addr),
    .R0_clk(mem_28_4_R0_clk),
    .R0_data(mem_28_4_R0_data),
    .R0_en(mem_28_4_R0_en),
    .W0_addr(mem_28_4_W0_addr),
    .W0_clk(mem_28_4_W0_clk),
    .W0_data(mem_28_4_W0_data),
    .W0_en(mem_28_4_W0_en),
    .W0_mask(mem_28_4_W0_mask)
  );
  split_mem_0_ext mem_28_5 (
    .R0_addr(mem_28_5_R0_addr),
    .R0_clk(mem_28_5_R0_clk),
    .R0_data(mem_28_5_R0_data),
    .R0_en(mem_28_5_R0_en),
    .W0_addr(mem_28_5_W0_addr),
    .W0_clk(mem_28_5_W0_clk),
    .W0_data(mem_28_5_W0_data),
    .W0_en(mem_28_5_W0_en),
    .W0_mask(mem_28_5_W0_mask)
  );
  split_mem_0_ext mem_28_6 (
    .R0_addr(mem_28_6_R0_addr),
    .R0_clk(mem_28_6_R0_clk),
    .R0_data(mem_28_6_R0_data),
    .R0_en(mem_28_6_R0_en),
    .W0_addr(mem_28_6_W0_addr),
    .W0_clk(mem_28_6_W0_clk),
    .W0_data(mem_28_6_W0_data),
    .W0_en(mem_28_6_W0_en),
    .W0_mask(mem_28_6_W0_mask)
  );
  split_mem_0_ext mem_28_7 (
    .R0_addr(mem_28_7_R0_addr),
    .R0_clk(mem_28_7_R0_clk),
    .R0_data(mem_28_7_R0_data),
    .R0_en(mem_28_7_R0_en),
    .W0_addr(mem_28_7_W0_addr),
    .W0_clk(mem_28_7_W0_clk),
    .W0_data(mem_28_7_W0_data),
    .W0_en(mem_28_7_W0_en),
    .W0_mask(mem_28_7_W0_mask)
  );
  split_mem_0_ext mem_29_0 (
    .R0_addr(mem_29_0_R0_addr),
    .R0_clk(mem_29_0_R0_clk),
    .R0_data(mem_29_0_R0_data),
    .R0_en(mem_29_0_R0_en),
    .W0_addr(mem_29_0_W0_addr),
    .W0_clk(mem_29_0_W0_clk),
    .W0_data(mem_29_0_W0_data),
    .W0_en(mem_29_0_W0_en),
    .W0_mask(mem_29_0_W0_mask)
  );
  split_mem_0_ext mem_29_1 (
    .R0_addr(mem_29_1_R0_addr),
    .R0_clk(mem_29_1_R0_clk),
    .R0_data(mem_29_1_R0_data),
    .R0_en(mem_29_1_R0_en),
    .W0_addr(mem_29_1_W0_addr),
    .W0_clk(mem_29_1_W0_clk),
    .W0_data(mem_29_1_W0_data),
    .W0_en(mem_29_1_W0_en),
    .W0_mask(mem_29_1_W0_mask)
  );
  split_mem_0_ext mem_29_2 (
    .R0_addr(mem_29_2_R0_addr),
    .R0_clk(mem_29_2_R0_clk),
    .R0_data(mem_29_2_R0_data),
    .R0_en(mem_29_2_R0_en),
    .W0_addr(mem_29_2_W0_addr),
    .W0_clk(mem_29_2_W0_clk),
    .W0_data(mem_29_2_W0_data),
    .W0_en(mem_29_2_W0_en),
    .W0_mask(mem_29_2_W0_mask)
  );
  split_mem_0_ext mem_29_3 (
    .R0_addr(mem_29_3_R0_addr),
    .R0_clk(mem_29_3_R0_clk),
    .R0_data(mem_29_3_R0_data),
    .R0_en(mem_29_3_R0_en),
    .W0_addr(mem_29_3_W0_addr),
    .W0_clk(mem_29_3_W0_clk),
    .W0_data(mem_29_3_W0_data),
    .W0_en(mem_29_3_W0_en),
    .W0_mask(mem_29_3_W0_mask)
  );
  split_mem_0_ext mem_29_4 (
    .R0_addr(mem_29_4_R0_addr),
    .R0_clk(mem_29_4_R0_clk),
    .R0_data(mem_29_4_R0_data),
    .R0_en(mem_29_4_R0_en),
    .W0_addr(mem_29_4_W0_addr),
    .W0_clk(mem_29_4_W0_clk),
    .W0_data(mem_29_4_W0_data),
    .W0_en(mem_29_4_W0_en),
    .W0_mask(mem_29_4_W0_mask)
  );
  split_mem_0_ext mem_29_5 (
    .R0_addr(mem_29_5_R0_addr),
    .R0_clk(mem_29_5_R0_clk),
    .R0_data(mem_29_5_R0_data),
    .R0_en(mem_29_5_R0_en),
    .W0_addr(mem_29_5_W0_addr),
    .W0_clk(mem_29_5_W0_clk),
    .W0_data(mem_29_5_W0_data),
    .W0_en(mem_29_5_W0_en),
    .W0_mask(mem_29_5_W0_mask)
  );
  split_mem_0_ext mem_29_6 (
    .R0_addr(mem_29_6_R0_addr),
    .R0_clk(mem_29_6_R0_clk),
    .R0_data(mem_29_6_R0_data),
    .R0_en(mem_29_6_R0_en),
    .W0_addr(mem_29_6_W0_addr),
    .W0_clk(mem_29_6_W0_clk),
    .W0_data(mem_29_6_W0_data),
    .W0_en(mem_29_6_W0_en),
    .W0_mask(mem_29_6_W0_mask)
  );
  split_mem_0_ext mem_29_7 (
    .R0_addr(mem_29_7_R0_addr),
    .R0_clk(mem_29_7_R0_clk),
    .R0_data(mem_29_7_R0_data),
    .R0_en(mem_29_7_R0_en),
    .W0_addr(mem_29_7_W0_addr),
    .W0_clk(mem_29_7_W0_clk),
    .W0_data(mem_29_7_W0_data),
    .W0_en(mem_29_7_W0_en),
    .W0_mask(mem_29_7_W0_mask)
  );
  split_mem_0_ext mem_30_0 (
    .R0_addr(mem_30_0_R0_addr),
    .R0_clk(mem_30_0_R0_clk),
    .R0_data(mem_30_0_R0_data),
    .R0_en(mem_30_0_R0_en),
    .W0_addr(mem_30_0_W0_addr),
    .W0_clk(mem_30_0_W0_clk),
    .W0_data(mem_30_0_W0_data),
    .W0_en(mem_30_0_W0_en),
    .W0_mask(mem_30_0_W0_mask)
  );
  split_mem_0_ext mem_30_1 (
    .R0_addr(mem_30_1_R0_addr),
    .R0_clk(mem_30_1_R0_clk),
    .R0_data(mem_30_1_R0_data),
    .R0_en(mem_30_1_R0_en),
    .W0_addr(mem_30_1_W0_addr),
    .W0_clk(mem_30_1_W0_clk),
    .W0_data(mem_30_1_W0_data),
    .W0_en(mem_30_1_W0_en),
    .W0_mask(mem_30_1_W0_mask)
  );
  split_mem_0_ext mem_30_2 (
    .R0_addr(mem_30_2_R0_addr),
    .R0_clk(mem_30_2_R0_clk),
    .R0_data(mem_30_2_R0_data),
    .R0_en(mem_30_2_R0_en),
    .W0_addr(mem_30_2_W0_addr),
    .W0_clk(mem_30_2_W0_clk),
    .W0_data(mem_30_2_W0_data),
    .W0_en(mem_30_2_W0_en),
    .W0_mask(mem_30_2_W0_mask)
  );
  split_mem_0_ext mem_30_3 (
    .R0_addr(mem_30_3_R0_addr),
    .R0_clk(mem_30_3_R0_clk),
    .R0_data(mem_30_3_R0_data),
    .R0_en(mem_30_3_R0_en),
    .W0_addr(mem_30_3_W0_addr),
    .W0_clk(mem_30_3_W0_clk),
    .W0_data(mem_30_3_W0_data),
    .W0_en(mem_30_3_W0_en),
    .W0_mask(mem_30_3_W0_mask)
  );
  split_mem_0_ext mem_30_4 (
    .R0_addr(mem_30_4_R0_addr),
    .R0_clk(mem_30_4_R0_clk),
    .R0_data(mem_30_4_R0_data),
    .R0_en(mem_30_4_R0_en),
    .W0_addr(mem_30_4_W0_addr),
    .W0_clk(mem_30_4_W0_clk),
    .W0_data(mem_30_4_W0_data),
    .W0_en(mem_30_4_W0_en),
    .W0_mask(mem_30_4_W0_mask)
  );
  split_mem_0_ext mem_30_5 (
    .R0_addr(mem_30_5_R0_addr),
    .R0_clk(mem_30_5_R0_clk),
    .R0_data(mem_30_5_R0_data),
    .R0_en(mem_30_5_R0_en),
    .W0_addr(mem_30_5_W0_addr),
    .W0_clk(mem_30_5_W0_clk),
    .W0_data(mem_30_5_W0_data),
    .W0_en(mem_30_5_W0_en),
    .W0_mask(mem_30_5_W0_mask)
  );
  split_mem_0_ext mem_30_6 (
    .R0_addr(mem_30_6_R0_addr),
    .R0_clk(mem_30_6_R0_clk),
    .R0_data(mem_30_6_R0_data),
    .R0_en(mem_30_6_R0_en),
    .W0_addr(mem_30_6_W0_addr),
    .W0_clk(mem_30_6_W0_clk),
    .W0_data(mem_30_6_W0_data),
    .W0_en(mem_30_6_W0_en),
    .W0_mask(mem_30_6_W0_mask)
  );
  split_mem_0_ext mem_30_7 (
    .R0_addr(mem_30_7_R0_addr),
    .R0_clk(mem_30_7_R0_clk),
    .R0_data(mem_30_7_R0_data),
    .R0_en(mem_30_7_R0_en),
    .W0_addr(mem_30_7_W0_addr),
    .W0_clk(mem_30_7_W0_clk),
    .W0_data(mem_30_7_W0_data),
    .W0_en(mem_30_7_W0_en),
    .W0_mask(mem_30_7_W0_mask)
  );
  split_mem_0_ext mem_31_0 (
    .R0_addr(mem_31_0_R0_addr),
    .R0_clk(mem_31_0_R0_clk),
    .R0_data(mem_31_0_R0_data),
    .R0_en(mem_31_0_R0_en),
    .W0_addr(mem_31_0_W0_addr),
    .W0_clk(mem_31_0_W0_clk),
    .W0_data(mem_31_0_W0_data),
    .W0_en(mem_31_0_W0_en),
    .W0_mask(mem_31_0_W0_mask)
  );
  split_mem_0_ext mem_31_1 (
    .R0_addr(mem_31_1_R0_addr),
    .R0_clk(mem_31_1_R0_clk),
    .R0_data(mem_31_1_R0_data),
    .R0_en(mem_31_1_R0_en),
    .W0_addr(mem_31_1_W0_addr),
    .W0_clk(mem_31_1_W0_clk),
    .W0_data(mem_31_1_W0_data),
    .W0_en(mem_31_1_W0_en),
    .W0_mask(mem_31_1_W0_mask)
  );
  split_mem_0_ext mem_31_2 (
    .R0_addr(mem_31_2_R0_addr),
    .R0_clk(mem_31_2_R0_clk),
    .R0_data(mem_31_2_R0_data),
    .R0_en(mem_31_2_R0_en),
    .W0_addr(mem_31_2_W0_addr),
    .W0_clk(mem_31_2_W0_clk),
    .W0_data(mem_31_2_W0_data),
    .W0_en(mem_31_2_W0_en),
    .W0_mask(mem_31_2_W0_mask)
  );
  split_mem_0_ext mem_31_3 (
    .R0_addr(mem_31_3_R0_addr),
    .R0_clk(mem_31_3_R0_clk),
    .R0_data(mem_31_3_R0_data),
    .R0_en(mem_31_3_R0_en),
    .W0_addr(mem_31_3_W0_addr),
    .W0_clk(mem_31_3_W0_clk),
    .W0_data(mem_31_3_W0_data),
    .W0_en(mem_31_3_W0_en),
    .W0_mask(mem_31_3_W0_mask)
  );
  split_mem_0_ext mem_31_4 (
    .R0_addr(mem_31_4_R0_addr),
    .R0_clk(mem_31_4_R0_clk),
    .R0_data(mem_31_4_R0_data),
    .R0_en(mem_31_4_R0_en),
    .W0_addr(mem_31_4_W0_addr),
    .W0_clk(mem_31_4_W0_clk),
    .W0_data(mem_31_4_W0_data),
    .W0_en(mem_31_4_W0_en),
    .W0_mask(mem_31_4_W0_mask)
  );
  split_mem_0_ext mem_31_5 (
    .R0_addr(mem_31_5_R0_addr),
    .R0_clk(mem_31_5_R0_clk),
    .R0_data(mem_31_5_R0_data),
    .R0_en(mem_31_5_R0_en),
    .W0_addr(mem_31_5_W0_addr),
    .W0_clk(mem_31_5_W0_clk),
    .W0_data(mem_31_5_W0_data),
    .W0_en(mem_31_5_W0_en),
    .W0_mask(mem_31_5_W0_mask)
  );
  split_mem_0_ext mem_31_6 (
    .R0_addr(mem_31_6_R0_addr),
    .R0_clk(mem_31_6_R0_clk),
    .R0_data(mem_31_6_R0_data),
    .R0_en(mem_31_6_R0_en),
    .W0_addr(mem_31_6_W0_addr),
    .W0_clk(mem_31_6_W0_clk),
    .W0_data(mem_31_6_W0_data),
    .W0_en(mem_31_6_W0_en),
    .W0_mask(mem_31_6_W0_mask)
  );
  split_mem_0_ext mem_31_7 (
    .R0_addr(mem_31_7_R0_addr),
    .R0_clk(mem_31_7_R0_clk),
    .R0_data(mem_31_7_R0_data),
    .R0_en(mem_31_7_R0_en),
    .W0_addr(mem_31_7_W0_addr),
    .W0_clk(mem_31_7_W0_clk),
    .W0_data(mem_31_7_W0_data),
    .W0_en(mem_31_7_W0_en),
    .W0_mask(mem_31_7_W0_mask)
  );
  split_mem_0_ext mem_32_0 (
    .R0_addr(mem_32_0_R0_addr),
    .R0_clk(mem_32_0_R0_clk),
    .R0_data(mem_32_0_R0_data),
    .R0_en(mem_32_0_R0_en),
    .W0_addr(mem_32_0_W0_addr),
    .W0_clk(mem_32_0_W0_clk),
    .W0_data(mem_32_0_W0_data),
    .W0_en(mem_32_0_W0_en),
    .W0_mask(mem_32_0_W0_mask)
  );
  split_mem_0_ext mem_32_1 (
    .R0_addr(mem_32_1_R0_addr),
    .R0_clk(mem_32_1_R0_clk),
    .R0_data(mem_32_1_R0_data),
    .R0_en(mem_32_1_R0_en),
    .W0_addr(mem_32_1_W0_addr),
    .W0_clk(mem_32_1_W0_clk),
    .W0_data(mem_32_1_W0_data),
    .W0_en(mem_32_1_W0_en),
    .W0_mask(mem_32_1_W0_mask)
  );
  split_mem_0_ext mem_32_2 (
    .R0_addr(mem_32_2_R0_addr),
    .R0_clk(mem_32_2_R0_clk),
    .R0_data(mem_32_2_R0_data),
    .R0_en(mem_32_2_R0_en),
    .W0_addr(mem_32_2_W0_addr),
    .W0_clk(mem_32_2_W0_clk),
    .W0_data(mem_32_2_W0_data),
    .W0_en(mem_32_2_W0_en),
    .W0_mask(mem_32_2_W0_mask)
  );
  split_mem_0_ext mem_32_3 (
    .R0_addr(mem_32_3_R0_addr),
    .R0_clk(mem_32_3_R0_clk),
    .R0_data(mem_32_3_R0_data),
    .R0_en(mem_32_3_R0_en),
    .W0_addr(mem_32_3_W0_addr),
    .W0_clk(mem_32_3_W0_clk),
    .W0_data(mem_32_3_W0_data),
    .W0_en(mem_32_3_W0_en),
    .W0_mask(mem_32_3_W0_mask)
  );
  split_mem_0_ext mem_32_4 (
    .R0_addr(mem_32_4_R0_addr),
    .R0_clk(mem_32_4_R0_clk),
    .R0_data(mem_32_4_R0_data),
    .R0_en(mem_32_4_R0_en),
    .W0_addr(mem_32_4_W0_addr),
    .W0_clk(mem_32_4_W0_clk),
    .W0_data(mem_32_4_W0_data),
    .W0_en(mem_32_4_W0_en),
    .W0_mask(mem_32_4_W0_mask)
  );
  split_mem_0_ext mem_32_5 (
    .R0_addr(mem_32_5_R0_addr),
    .R0_clk(mem_32_5_R0_clk),
    .R0_data(mem_32_5_R0_data),
    .R0_en(mem_32_5_R0_en),
    .W0_addr(mem_32_5_W0_addr),
    .W0_clk(mem_32_5_W0_clk),
    .W0_data(mem_32_5_W0_data),
    .W0_en(mem_32_5_W0_en),
    .W0_mask(mem_32_5_W0_mask)
  );
  split_mem_0_ext mem_32_6 (
    .R0_addr(mem_32_6_R0_addr),
    .R0_clk(mem_32_6_R0_clk),
    .R0_data(mem_32_6_R0_data),
    .R0_en(mem_32_6_R0_en),
    .W0_addr(mem_32_6_W0_addr),
    .W0_clk(mem_32_6_W0_clk),
    .W0_data(mem_32_6_W0_data),
    .W0_en(mem_32_6_W0_en),
    .W0_mask(mem_32_6_W0_mask)
  );
  split_mem_0_ext mem_32_7 (
    .R0_addr(mem_32_7_R0_addr),
    .R0_clk(mem_32_7_R0_clk),
    .R0_data(mem_32_7_R0_data),
    .R0_en(mem_32_7_R0_en),
    .W0_addr(mem_32_7_W0_addr),
    .W0_clk(mem_32_7_W0_clk),
    .W0_data(mem_32_7_W0_data),
    .W0_en(mem_32_7_W0_en),
    .W0_mask(mem_32_7_W0_mask)
  );
  split_mem_0_ext mem_33_0 (
    .R0_addr(mem_33_0_R0_addr),
    .R0_clk(mem_33_0_R0_clk),
    .R0_data(mem_33_0_R0_data),
    .R0_en(mem_33_0_R0_en),
    .W0_addr(mem_33_0_W0_addr),
    .W0_clk(mem_33_0_W0_clk),
    .W0_data(mem_33_0_W0_data),
    .W0_en(mem_33_0_W0_en),
    .W0_mask(mem_33_0_W0_mask)
  );
  split_mem_0_ext mem_33_1 (
    .R0_addr(mem_33_1_R0_addr),
    .R0_clk(mem_33_1_R0_clk),
    .R0_data(mem_33_1_R0_data),
    .R0_en(mem_33_1_R0_en),
    .W0_addr(mem_33_1_W0_addr),
    .W0_clk(mem_33_1_W0_clk),
    .W0_data(mem_33_1_W0_data),
    .W0_en(mem_33_1_W0_en),
    .W0_mask(mem_33_1_W0_mask)
  );
  split_mem_0_ext mem_33_2 (
    .R0_addr(mem_33_2_R0_addr),
    .R0_clk(mem_33_2_R0_clk),
    .R0_data(mem_33_2_R0_data),
    .R0_en(mem_33_2_R0_en),
    .W0_addr(mem_33_2_W0_addr),
    .W0_clk(mem_33_2_W0_clk),
    .W0_data(mem_33_2_W0_data),
    .W0_en(mem_33_2_W0_en),
    .W0_mask(mem_33_2_W0_mask)
  );
  split_mem_0_ext mem_33_3 (
    .R0_addr(mem_33_3_R0_addr),
    .R0_clk(mem_33_3_R0_clk),
    .R0_data(mem_33_3_R0_data),
    .R0_en(mem_33_3_R0_en),
    .W0_addr(mem_33_3_W0_addr),
    .W0_clk(mem_33_3_W0_clk),
    .W0_data(mem_33_3_W0_data),
    .W0_en(mem_33_3_W0_en),
    .W0_mask(mem_33_3_W0_mask)
  );
  split_mem_0_ext mem_33_4 (
    .R0_addr(mem_33_4_R0_addr),
    .R0_clk(mem_33_4_R0_clk),
    .R0_data(mem_33_4_R0_data),
    .R0_en(mem_33_4_R0_en),
    .W0_addr(mem_33_4_W0_addr),
    .W0_clk(mem_33_4_W0_clk),
    .W0_data(mem_33_4_W0_data),
    .W0_en(mem_33_4_W0_en),
    .W0_mask(mem_33_4_W0_mask)
  );
  split_mem_0_ext mem_33_5 (
    .R0_addr(mem_33_5_R0_addr),
    .R0_clk(mem_33_5_R0_clk),
    .R0_data(mem_33_5_R0_data),
    .R0_en(mem_33_5_R0_en),
    .W0_addr(mem_33_5_W0_addr),
    .W0_clk(mem_33_5_W0_clk),
    .W0_data(mem_33_5_W0_data),
    .W0_en(mem_33_5_W0_en),
    .W0_mask(mem_33_5_W0_mask)
  );
  split_mem_0_ext mem_33_6 (
    .R0_addr(mem_33_6_R0_addr),
    .R0_clk(mem_33_6_R0_clk),
    .R0_data(mem_33_6_R0_data),
    .R0_en(mem_33_6_R0_en),
    .W0_addr(mem_33_6_W0_addr),
    .W0_clk(mem_33_6_W0_clk),
    .W0_data(mem_33_6_W0_data),
    .W0_en(mem_33_6_W0_en),
    .W0_mask(mem_33_6_W0_mask)
  );
  split_mem_0_ext mem_33_7 (
    .R0_addr(mem_33_7_R0_addr),
    .R0_clk(mem_33_7_R0_clk),
    .R0_data(mem_33_7_R0_data),
    .R0_en(mem_33_7_R0_en),
    .W0_addr(mem_33_7_W0_addr),
    .W0_clk(mem_33_7_W0_clk),
    .W0_data(mem_33_7_W0_data),
    .W0_en(mem_33_7_W0_en),
    .W0_mask(mem_33_7_W0_mask)
  );
  split_mem_0_ext mem_34_0 (
    .R0_addr(mem_34_0_R0_addr),
    .R0_clk(mem_34_0_R0_clk),
    .R0_data(mem_34_0_R0_data),
    .R0_en(mem_34_0_R0_en),
    .W0_addr(mem_34_0_W0_addr),
    .W0_clk(mem_34_0_W0_clk),
    .W0_data(mem_34_0_W0_data),
    .W0_en(mem_34_0_W0_en),
    .W0_mask(mem_34_0_W0_mask)
  );
  split_mem_0_ext mem_34_1 (
    .R0_addr(mem_34_1_R0_addr),
    .R0_clk(mem_34_1_R0_clk),
    .R0_data(mem_34_1_R0_data),
    .R0_en(mem_34_1_R0_en),
    .W0_addr(mem_34_1_W0_addr),
    .W0_clk(mem_34_1_W0_clk),
    .W0_data(mem_34_1_W0_data),
    .W0_en(mem_34_1_W0_en),
    .W0_mask(mem_34_1_W0_mask)
  );
  split_mem_0_ext mem_34_2 (
    .R0_addr(mem_34_2_R0_addr),
    .R0_clk(mem_34_2_R0_clk),
    .R0_data(mem_34_2_R0_data),
    .R0_en(mem_34_2_R0_en),
    .W0_addr(mem_34_2_W0_addr),
    .W0_clk(mem_34_2_W0_clk),
    .W0_data(mem_34_2_W0_data),
    .W0_en(mem_34_2_W0_en),
    .W0_mask(mem_34_2_W0_mask)
  );
  split_mem_0_ext mem_34_3 (
    .R0_addr(mem_34_3_R0_addr),
    .R0_clk(mem_34_3_R0_clk),
    .R0_data(mem_34_3_R0_data),
    .R0_en(mem_34_3_R0_en),
    .W0_addr(mem_34_3_W0_addr),
    .W0_clk(mem_34_3_W0_clk),
    .W0_data(mem_34_3_W0_data),
    .W0_en(mem_34_3_W0_en),
    .W0_mask(mem_34_3_W0_mask)
  );
  split_mem_0_ext mem_34_4 (
    .R0_addr(mem_34_4_R0_addr),
    .R0_clk(mem_34_4_R0_clk),
    .R0_data(mem_34_4_R0_data),
    .R0_en(mem_34_4_R0_en),
    .W0_addr(mem_34_4_W0_addr),
    .W0_clk(mem_34_4_W0_clk),
    .W0_data(mem_34_4_W0_data),
    .W0_en(mem_34_4_W0_en),
    .W0_mask(mem_34_4_W0_mask)
  );
  split_mem_0_ext mem_34_5 (
    .R0_addr(mem_34_5_R0_addr),
    .R0_clk(mem_34_5_R0_clk),
    .R0_data(mem_34_5_R0_data),
    .R0_en(mem_34_5_R0_en),
    .W0_addr(mem_34_5_W0_addr),
    .W0_clk(mem_34_5_W0_clk),
    .W0_data(mem_34_5_W0_data),
    .W0_en(mem_34_5_W0_en),
    .W0_mask(mem_34_5_W0_mask)
  );
  split_mem_0_ext mem_34_6 (
    .R0_addr(mem_34_6_R0_addr),
    .R0_clk(mem_34_6_R0_clk),
    .R0_data(mem_34_6_R0_data),
    .R0_en(mem_34_6_R0_en),
    .W0_addr(mem_34_6_W0_addr),
    .W0_clk(mem_34_6_W0_clk),
    .W0_data(mem_34_6_W0_data),
    .W0_en(mem_34_6_W0_en),
    .W0_mask(mem_34_6_W0_mask)
  );
  split_mem_0_ext mem_34_7 (
    .R0_addr(mem_34_7_R0_addr),
    .R0_clk(mem_34_7_R0_clk),
    .R0_data(mem_34_7_R0_data),
    .R0_en(mem_34_7_R0_en),
    .W0_addr(mem_34_7_W0_addr),
    .W0_clk(mem_34_7_W0_clk),
    .W0_data(mem_34_7_W0_data),
    .W0_en(mem_34_7_W0_en),
    .W0_mask(mem_34_7_W0_mask)
  );
  split_mem_0_ext mem_35_0 (
    .R0_addr(mem_35_0_R0_addr),
    .R0_clk(mem_35_0_R0_clk),
    .R0_data(mem_35_0_R0_data),
    .R0_en(mem_35_0_R0_en),
    .W0_addr(mem_35_0_W0_addr),
    .W0_clk(mem_35_0_W0_clk),
    .W0_data(mem_35_0_W0_data),
    .W0_en(mem_35_0_W0_en),
    .W0_mask(mem_35_0_W0_mask)
  );
  split_mem_0_ext mem_35_1 (
    .R0_addr(mem_35_1_R0_addr),
    .R0_clk(mem_35_1_R0_clk),
    .R0_data(mem_35_1_R0_data),
    .R0_en(mem_35_1_R0_en),
    .W0_addr(mem_35_1_W0_addr),
    .W0_clk(mem_35_1_W0_clk),
    .W0_data(mem_35_1_W0_data),
    .W0_en(mem_35_1_W0_en),
    .W0_mask(mem_35_1_W0_mask)
  );
  split_mem_0_ext mem_35_2 (
    .R0_addr(mem_35_2_R0_addr),
    .R0_clk(mem_35_2_R0_clk),
    .R0_data(mem_35_2_R0_data),
    .R0_en(mem_35_2_R0_en),
    .W0_addr(mem_35_2_W0_addr),
    .W0_clk(mem_35_2_W0_clk),
    .W0_data(mem_35_2_W0_data),
    .W0_en(mem_35_2_W0_en),
    .W0_mask(mem_35_2_W0_mask)
  );
  split_mem_0_ext mem_35_3 (
    .R0_addr(mem_35_3_R0_addr),
    .R0_clk(mem_35_3_R0_clk),
    .R0_data(mem_35_3_R0_data),
    .R0_en(mem_35_3_R0_en),
    .W0_addr(mem_35_3_W0_addr),
    .W0_clk(mem_35_3_W0_clk),
    .W0_data(mem_35_3_W0_data),
    .W0_en(mem_35_3_W0_en),
    .W0_mask(mem_35_3_W0_mask)
  );
  split_mem_0_ext mem_35_4 (
    .R0_addr(mem_35_4_R0_addr),
    .R0_clk(mem_35_4_R0_clk),
    .R0_data(mem_35_4_R0_data),
    .R0_en(mem_35_4_R0_en),
    .W0_addr(mem_35_4_W0_addr),
    .W0_clk(mem_35_4_W0_clk),
    .W0_data(mem_35_4_W0_data),
    .W0_en(mem_35_4_W0_en),
    .W0_mask(mem_35_4_W0_mask)
  );
  split_mem_0_ext mem_35_5 (
    .R0_addr(mem_35_5_R0_addr),
    .R0_clk(mem_35_5_R0_clk),
    .R0_data(mem_35_5_R0_data),
    .R0_en(mem_35_5_R0_en),
    .W0_addr(mem_35_5_W0_addr),
    .W0_clk(mem_35_5_W0_clk),
    .W0_data(mem_35_5_W0_data),
    .W0_en(mem_35_5_W0_en),
    .W0_mask(mem_35_5_W0_mask)
  );
  split_mem_0_ext mem_35_6 (
    .R0_addr(mem_35_6_R0_addr),
    .R0_clk(mem_35_6_R0_clk),
    .R0_data(mem_35_6_R0_data),
    .R0_en(mem_35_6_R0_en),
    .W0_addr(mem_35_6_W0_addr),
    .W0_clk(mem_35_6_W0_clk),
    .W0_data(mem_35_6_W0_data),
    .W0_en(mem_35_6_W0_en),
    .W0_mask(mem_35_6_W0_mask)
  );
  split_mem_0_ext mem_35_7 (
    .R0_addr(mem_35_7_R0_addr),
    .R0_clk(mem_35_7_R0_clk),
    .R0_data(mem_35_7_R0_data),
    .R0_en(mem_35_7_R0_en),
    .W0_addr(mem_35_7_W0_addr),
    .W0_clk(mem_35_7_W0_clk),
    .W0_data(mem_35_7_W0_data),
    .W0_en(mem_35_7_W0_en),
    .W0_mask(mem_35_7_W0_mask)
  );
  split_mem_0_ext mem_36_0 (
    .R0_addr(mem_36_0_R0_addr),
    .R0_clk(mem_36_0_R0_clk),
    .R0_data(mem_36_0_R0_data),
    .R0_en(mem_36_0_R0_en),
    .W0_addr(mem_36_0_W0_addr),
    .W0_clk(mem_36_0_W0_clk),
    .W0_data(mem_36_0_W0_data),
    .W0_en(mem_36_0_W0_en),
    .W0_mask(mem_36_0_W0_mask)
  );
  split_mem_0_ext mem_36_1 (
    .R0_addr(mem_36_1_R0_addr),
    .R0_clk(mem_36_1_R0_clk),
    .R0_data(mem_36_1_R0_data),
    .R0_en(mem_36_1_R0_en),
    .W0_addr(mem_36_1_W0_addr),
    .W0_clk(mem_36_1_W0_clk),
    .W0_data(mem_36_1_W0_data),
    .W0_en(mem_36_1_W0_en),
    .W0_mask(mem_36_1_W0_mask)
  );
  split_mem_0_ext mem_36_2 (
    .R0_addr(mem_36_2_R0_addr),
    .R0_clk(mem_36_2_R0_clk),
    .R0_data(mem_36_2_R0_data),
    .R0_en(mem_36_2_R0_en),
    .W0_addr(mem_36_2_W0_addr),
    .W0_clk(mem_36_2_W0_clk),
    .W0_data(mem_36_2_W0_data),
    .W0_en(mem_36_2_W0_en),
    .W0_mask(mem_36_2_W0_mask)
  );
  split_mem_0_ext mem_36_3 (
    .R0_addr(mem_36_3_R0_addr),
    .R0_clk(mem_36_3_R0_clk),
    .R0_data(mem_36_3_R0_data),
    .R0_en(mem_36_3_R0_en),
    .W0_addr(mem_36_3_W0_addr),
    .W0_clk(mem_36_3_W0_clk),
    .W0_data(mem_36_3_W0_data),
    .W0_en(mem_36_3_W0_en),
    .W0_mask(mem_36_3_W0_mask)
  );
  split_mem_0_ext mem_36_4 (
    .R0_addr(mem_36_4_R0_addr),
    .R0_clk(mem_36_4_R0_clk),
    .R0_data(mem_36_4_R0_data),
    .R0_en(mem_36_4_R0_en),
    .W0_addr(mem_36_4_W0_addr),
    .W0_clk(mem_36_4_W0_clk),
    .W0_data(mem_36_4_W0_data),
    .W0_en(mem_36_4_W0_en),
    .W0_mask(mem_36_4_W0_mask)
  );
  split_mem_0_ext mem_36_5 (
    .R0_addr(mem_36_5_R0_addr),
    .R0_clk(mem_36_5_R0_clk),
    .R0_data(mem_36_5_R0_data),
    .R0_en(mem_36_5_R0_en),
    .W0_addr(mem_36_5_W0_addr),
    .W0_clk(mem_36_5_W0_clk),
    .W0_data(mem_36_5_W0_data),
    .W0_en(mem_36_5_W0_en),
    .W0_mask(mem_36_5_W0_mask)
  );
  split_mem_0_ext mem_36_6 (
    .R0_addr(mem_36_6_R0_addr),
    .R0_clk(mem_36_6_R0_clk),
    .R0_data(mem_36_6_R0_data),
    .R0_en(mem_36_6_R0_en),
    .W0_addr(mem_36_6_W0_addr),
    .W0_clk(mem_36_6_W0_clk),
    .W0_data(mem_36_6_W0_data),
    .W0_en(mem_36_6_W0_en),
    .W0_mask(mem_36_6_W0_mask)
  );
  split_mem_0_ext mem_36_7 (
    .R0_addr(mem_36_7_R0_addr),
    .R0_clk(mem_36_7_R0_clk),
    .R0_data(mem_36_7_R0_data),
    .R0_en(mem_36_7_R0_en),
    .W0_addr(mem_36_7_W0_addr),
    .W0_clk(mem_36_7_W0_clk),
    .W0_data(mem_36_7_W0_data),
    .W0_en(mem_36_7_W0_en),
    .W0_mask(mem_36_7_W0_mask)
  );
  split_mem_0_ext mem_37_0 (
    .R0_addr(mem_37_0_R0_addr),
    .R0_clk(mem_37_0_R0_clk),
    .R0_data(mem_37_0_R0_data),
    .R0_en(mem_37_0_R0_en),
    .W0_addr(mem_37_0_W0_addr),
    .W0_clk(mem_37_0_W0_clk),
    .W0_data(mem_37_0_W0_data),
    .W0_en(mem_37_0_W0_en),
    .W0_mask(mem_37_0_W0_mask)
  );
  split_mem_0_ext mem_37_1 (
    .R0_addr(mem_37_1_R0_addr),
    .R0_clk(mem_37_1_R0_clk),
    .R0_data(mem_37_1_R0_data),
    .R0_en(mem_37_1_R0_en),
    .W0_addr(mem_37_1_W0_addr),
    .W0_clk(mem_37_1_W0_clk),
    .W0_data(mem_37_1_W0_data),
    .W0_en(mem_37_1_W0_en),
    .W0_mask(mem_37_1_W0_mask)
  );
  split_mem_0_ext mem_37_2 (
    .R0_addr(mem_37_2_R0_addr),
    .R0_clk(mem_37_2_R0_clk),
    .R0_data(mem_37_2_R0_data),
    .R0_en(mem_37_2_R0_en),
    .W0_addr(mem_37_2_W0_addr),
    .W0_clk(mem_37_2_W0_clk),
    .W0_data(mem_37_2_W0_data),
    .W0_en(mem_37_2_W0_en),
    .W0_mask(mem_37_2_W0_mask)
  );
  split_mem_0_ext mem_37_3 (
    .R0_addr(mem_37_3_R0_addr),
    .R0_clk(mem_37_3_R0_clk),
    .R0_data(mem_37_3_R0_data),
    .R0_en(mem_37_3_R0_en),
    .W0_addr(mem_37_3_W0_addr),
    .W0_clk(mem_37_3_W0_clk),
    .W0_data(mem_37_3_W0_data),
    .W0_en(mem_37_3_W0_en),
    .W0_mask(mem_37_3_W0_mask)
  );
  split_mem_0_ext mem_37_4 (
    .R0_addr(mem_37_4_R0_addr),
    .R0_clk(mem_37_4_R0_clk),
    .R0_data(mem_37_4_R0_data),
    .R0_en(mem_37_4_R0_en),
    .W0_addr(mem_37_4_W0_addr),
    .W0_clk(mem_37_4_W0_clk),
    .W0_data(mem_37_4_W0_data),
    .W0_en(mem_37_4_W0_en),
    .W0_mask(mem_37_4_W0_mask)
  );
  split_mem_0_ext mem_37_5 (
    .R0_addr(mem_37_5_R0_addr),
    .R0_clk(mem_37_5_R0_clk),
    .R0_data(mem_37_5_R0_data),
    .R0_en(mem_37_5_R0_en),
    .W0_addr(mem_37_5_W0_addr),
    .W0_clk(mem_37_5_W0_clk),
    .W0_data(mem_37_5_W0_data),
    .W0_en(mem_37_5_W0_en),
    .W0_mask(mem_37_5_W0_mask)
  );
  split_mem_0_ext mem_37_6 (
    .R0_addr(mem_37_6_R0_addr),
    .R0_clk(mem_37_6_R0_clk),
    .R0_data(mem_37_6_R0_data),
    .R0_en(mem_37_6_R0_en),
    .W0_addr(mem_37_6_W0_addr),
    .W0_clk(mem_37_6_W0_clk),
    .W0_data(mem_37_6_W0_data),
    .W0_en(mem_37_6_W0_en),
    .W0_mask(mem_37_6_W0_mask)
  );
  split_mem_0_ext mem_37_7 (
    .R0_addr(mem_37_7_R0_addr),
    .R0_clk(mem_37_7_R0_clk),
    .R0_data(mem_37_7_R0_data),
    .R0_en(mem_37_7_R0_en),
    .W0_addr(mem_37_7_W0_addr),
    .W0_clk(mem_37_7_W0_clk),
    .W0_data(mem_37_7_W0_data),
    .W0_en(mem_37_7_W0_en),
    .W0_mask(mem_37_7_W0_mask)
  );
  split_mem_0_ext mem_38_0 (
    .R0_addr(mem_38_0_R0_addr),
    .R0_clk(mem_38_0_R0_clk),
    .R0_data(mem_38_0_R0_data),
    .R0_en(mem_38_0_R0_en),
    .W0_addr(mem_38_0_W0_addr),
    .W0_clk(mem_38_0_W0_clk),
    .W0_data(mem_38_0_W0_data),
    .W0_en(mem_38_0_W0_en),
    .W0_mask(mem_38_0_W0_mask)
  );
  split_mem_0_ext mem_38_1 (
    .R0_addr(mem_38_1_R0_addr),
    .R0_clk(mem_38_1_R0_clk),
    .R0_data(mem_38_1_R0_data),
    .R0_en(mem_38_1_R0_en),
    .W0_addr(mem_38_1_W0_addr),
    .W0_clk(mem_38_1_W0_clk),
    .W0_data(mem_38_1_W0_data),
    .W0_en(mem_38_1_W0_en),
    .W0_mask(mem_38_1_W0_mask)
  );
  split_mem_0_ext mem_38_2 (
    .R0_addr(mem_38_2_R0_addr),
    .R0_clk(mem_38_2_R0_clk),
    .R0_data(mem_38_2_R0_data),
    .R0_en(mem_38_2_R0_en),
    .W0_addr(mem_38_2_W0_addr),
    .W0_clk(mem_38_2_W0_clk),
    .W0_data(mem_38_2_W0_data),
    .W0_en(mem_38_2_W0_en),
    .W0_mask(mem_38_2_W0_mask)
  );
  split_mem_0_ext mem_38_3 (
    .R0_addr(mem_38_3_R0_addr),
    .R0_clk(mem_38_3_R0_clk),
    .R0_data(mem_38_3_R0_data),
    .R0_en(mem_38_3_R0_en),
    .W0_addr(mem_38_3_W0_addr),
    .W0_clk(mem_38_3_W0_clk),
    .W0_data(mem_38_3_W0_data),
    .W0_en(mem_38_3_W0_en),
    .W0_mask(mem_38_3_W0_mask)
  );
  split_mem_0_ext mem_38_4 (
    .R0_addr(mem_38_4_R0_addr),
    .R0_clk(mem_38_4_R0_clk),
    .R0_data(mem_38_4_R0_data),
    .R0_en(mem_38_4_R0_en),
    .W0_addr(mem_38_4_W0_addr),
    .W0_clk(mem_38_4_W0_clk),
    .W0_data(mem_38_4_W0_data),
    .W0_en(mem_38_4_W0_en),
    .W0_mask(mem_38_4_W0_mask)
  );
  split_mem_0_ext mem_38_5 (
    .R0_addr(mem_38_5_R0_addr),
    .R0_clk(mem_38_5_R0_clk),
    .R0_data(mem_38_5_R0_data),
    .R0_en(mem_38_5_R0_en),
    .W0_addr(mem_38_5_W0_addr),
    .W0_clk(mem_38_5_W0_clk),
    .W0_data(mem_38_5_W0_data),
    .W0_en(mem_38_5_W0_en),
    .W0_mask(mem_38_5_W0_mask)
  );
  split_mem_0_ext mem_38_6 (
    .R0_addr(mem_38_6_R0_addr),
    .R0_clk(mem_38_6_R0_clk),
    .R0_data(mem_38_6_R0_data),
    .R0_en(mem_38_6_R0_en),
    .W0_addr(mem_38_6_W0_addr),
    .W0_clk(mem_38_6_W0_clk),
    .W0_data(mem_38_6_W0_data),
    .W0_en(mem_38_6_W0_en),
    .W0_mask(mem_38_6_W0_mask)
  );
  split_mem_0_ext mem_38_7 (
    .R0_addr(mem_38_7_R0_addr),
    .R0_clk(mem_38_7_R0_clk),
    .R0_data(mem_38_7_R0_data),
    .R0_en(mem_38_7_R0_en),
    .W0_addr(mem_38_7_W0_addr),
    .W0_clk(mem_38_7_W0_clk),
    .W0_data(mem_38_7_W0_data),
    .W0_en(mem_38_7_W0_en),
    .W0_mask(mem_38_7_W0_mask)
  );
  split_mem_0_ext mem_39_0 (
    .R0_addr(mem_39_0_R0_addr),
    .R0_clk(mem_39_0_R0_clk),
    .R0_data(mem_39_0_R0_data),
    .R0_en(mem_39_0_R0_en),
    .W0_addr(mem_39_0_W0_addr),
    .W0_clk(mem_39_0_W0_clk),
    .W0_data(mem_39_0_W0_data),
    .W0_en(mem_39_0_W0_en),
    .W0_mask(mem_39_0_W0_mask)
  );
  split_mem_0_ext mem_39_1 (
    .R0_addr(mem_39_1_R0_addr),
    .R0_clk(mem_39_1_R0_clk),
    .R0_data(mem_39_1_R0_data),
    .R0_en(mem_39_1_R0_en),
    .W0_addr(mem_39_1_W0_addr),
    .W0_clk(mem_39_1_W0_clk),
    .W0_data(mem_39_1_W0_data),
    .W0_en(mem_39_1_W0_en),
    .W0_mask(mem_39_1_W0_mask)
  );
  split_mem_0_ext mem_39_2 (
    .R0_addr(mem_39_2_R0_addr),
    .R0_clk(mem_39_2_R0_clk),
    .R0_data(mem_39_2_R0_data),
    .R0_en(mem_39_2_R0_en),
    .W0_addr(mem_39_2_W0_addr),
    .W0_clk(mem_39_2_W0_clk),
    .W0_data(mem_39_2_W0_data),
    .W0_en(mem_39_2_W0_en),
    .W0_mask(mem_39_2_W0_mask)
  );
  split_mem_0_ext mem_39_3 (
    .R0_addr(mem_39_3_R0_addr),
    .R0_clk(mem_39_3_R0_clk),
    .R0_data(mem_39_3_R0_data),
    .R0_en(mem_39_3_R0_en),
    .W0_addr(mem_39_3_W0_addr),
    .W0_clk(mem_39_3_W0_clk),
    .W0_data(mem_39_3_W0_data),
    .W0_en(mem_39_3_W0_en),
    .W0_mask(mem_39_3_W0_mask)
  );
  split_mem_0_ext mem_39_4 (
    .R0_addr(mem_39_4_R0_addr),
    .R0_clk(mem_39_4_R0_clk),
    .R0_data(mem_39_4_R0_data),
    .R0_en(mem_39_4_R0_en),
    .W0_addr(mem_39_4_W0_addr),
    .W0_clk(mem_39_4_W0_clk),
    .W0_data(mem_39_4_W0_data),
    .W0_en(mem_39_4_W0_en),
    .W0_mask(mem_39_4_W0_mask)
  );
  split_mem_0_ext mem_39_5 (
    .R0_addr(mem_39_5_R0_addr),
    .R0_clk(mem_39_5_R0_clk),
    .R0_data(mem_39_5_R0_data),
    .R0_en(mem_39_5_R0_en),
    .W0_addr(mem_39_5_W0_addr),
    .W0_clk(mem_39_5_W0_clk),
    .W0_data(mem_39_5_W0_data),
    .W0_en(mem_39_5_W0_en),
    .W0_mask(mem_39_5_W0_mask)
  );
  split_mem_0_ext mem_39_6 (
    .R0_addr(mem_39_6_R0_addr),
    .R0_clk(mem_39_6_R0_clk),
    .R0_data(mem_39_6_R0_data),
    .R0_en(mem_39_6_R0_en),
    .W0_addr(mem_39_6_W0_addr),
    .W0_clk(mem_39_6_W0_clk),
    .W0_data(mem_39_6_W0_data),
    .W0_en(mem_39_6_W0_en),
    .W0_mask(mem_39_6_W0_mask)
  );
  split_mem_0_ext mem_39_7 (
    .R0_addr(mem_39_7_R0_addr),
    .R0_clk(mem_39_7_R0_clk),
    .R0_data(mem_39_7_R0_data),
    .R0_en(mem_39_7_R0_en),
    .W0_addr(mem_39_7_W0_addr),
    .W0_clk(mem_39_7_W0_clk),
    .W0_data(mem_39_7_W0_data),
    .W0_en(mem_39_7_W0_en),
    .W0_mask(mem_39_7_W0_mask)
  );
  split_mem_0_ext mem_40_0 (
    .R0_addr(mem_40_0_R0_addr),
    .R0_clk(mem_40_0_R0_clk),
    .R0_data(mem_40_0_R0_data),
    .R0_en(mem_40_0_R0_en),
    .W0_addr(mem_40_0_W0_addr),
    .W0_clk(mem_40_0_W0_clk),
    .W0_data(mem_40_0_W0_data),
    .W0_en(mem_40_0_W0_en),
    .W0_mask(mem_40_0_W0_mask)
  );
  split_mem_0_ext mem_40_1 (
    .R0_addr(mem_40_1_R0_addr),
    .R0_clk(mem_40_1_R0_clk),
    .R0_data(mem_40_1_R0_data),
    .R0_en(mem_40_1_R0_en),
    .W0_addr(mem_40_1_W0_addr),
    .W0_clk(mem_40_1_W0_clk),
    .W0_data(mem_40_1_W0_data),
    .W0_en(mem_40_1_W0_en),
    .W0_mask(mem_40_1_W0_mask)
  );
  split_mem_0_ext mem_40_2 (
    .R0_addr(mem_40_2_R0_addr),
    .R0_clk(mem_40_2_R0_clk),
    .R0_data(mem_40_2_R0_data),
    .R0_en(mem_40_2_R0_en),
    .W0_addr(mem_40_2_W0_addr),
    .W0_clk(mem_40_2_W0_clk),
    .W0_data(mem_40_2_W0_data),
    .W0_en(mem_40_2_W0_en),
    .W0_mask(mem_40_2_W0_mask)
  );
  split_mem_0_ext mem_40_3 (
    .R0_addr(mem_40_3_R0_addr),
    .R0_clk(mem_40_3_R0_clk),
    .R0_data(mem_40_3_R0_data),
    .R0_en(mem_40_3_R0_en),
    .W0_addr(mem_40_3_W0_addr),
    .W0_clk(mem_40_3_W0_clk),
    .W0_data(mem_40_3_W0_data),
    .W0_en(mem_40_3_W0_en),
    .W0_mask(mem_40_3_W0_mask)
  );
  split_mem_0_ext mem_40_4 (
    .R0_addr(mem_40_4_R0_addr),
    .R0_clk(mem_40_4_R0_clk),
    .R0_data(mem_40_4_R0_data),
    .R0_en(mem_40_4_R0_en),
    .W0_addr(mem_40_4_W0_addr),
    .W0_clk(mem_40_4_W0_clk),
    .W0_data(mem_40_4_W0_data),
    .W0_en(mem_40_4_W0_en),
    .W0_mask(mem_40_4_W0_mask)
  );
  split_mem_0_ext mem_40_5 (
    .R0_addr(mem_40_5_R0_addr),
    .R0_clk(mem_40_5_R0_clk),
    .R0_data(mem_40_5_R0_data),
    .R0_en(mem_40_5_R0_en),
    .W0_addr(mem_40_5_W0_addr),
    .W0_clk(mem_40_5_W0_clk),
    .W0_data(mem_40_5_W0_data),
    .W0_en(mem_40_5_W0_en),
    .W0_mask(mem_40_5_W0_mask)
  );
  split_mem_0_ext mem_40_6 (
    .R0_addr(mem_40_6_R0_addr),
    .R0_clk(mem_40_6_R0_clk),
    .R0_data(mem_40_6_R0_data),
    .R0_en(mem_40_6_R0_en),
    .W0_addr(mem_40_6_W0_addr),
    .W0_clk(mem_40_6_W0_clk),
    .W0_data(mem_40_6_W0_data),
    .W0_en(mem_40_6_W0_en),
    .W0_mask(mem_40_6_W0_mask)
  );
  split_mem_0_ext mem_40_7 (
    .R0_addr(mem_40_7_R0_addr),
    .R0_clk(mem_40_7_R0_clk),
    .R0_data(mem_40_7_R0_data),
    .R0_en(mem_40_7_R0_en),
    .W0_addr(mem_40_7_W0_addr),
    .W0_clk(mem_40_7_W0_clk),
    .W0_data(mem_40_7_W0_data),
    .W0_en(mem_40_7_W0_en),
    .W0_mask(mem_40_7_W0_mask)
  );
  split_mem_0_ext mem_41_0 (
    .R0_addr(mem_41_0_R0_addr),
    .R0_clk(mem_41_0_R0_clk),
    .R0_data(mem_41_0_R0_data),
    .R0_en(mem_41_0_R0_en),
    .W0_addr(mem_41_0_W0_addr),
    .W0_clk(mem_41_0_W0_clk),
    .W0_data(mem_41_0_W0_data),
    .W0_en(mem_41_0_W0_en),
    .W0_mask(mem_41_0_W0_mask)
  );
  split_mem_0_ext mem_41_1 (
    .R0_addr(mem_41_1_R0_addr),
    .R0_clk(mem_41_1_R0_clk),
    .R0_data(mem_41_1_R0_data),
    .R0_en(mem_41_1_R0_en),
    .W0_addr(mem_41_1_W0_addr),
    .W0_clk(mem_41_1_W0_clk),
    .W0_data(mem_41_1_W0_data),
    .W0_en(mem_41_1_W0_en),
    .W0_mask(mem_41_1_W0_mask)
  );
  split_mem_0_ext mem_41_2 (
    .R0_addr(mem_41_2_R0_addr),
    .R0_clk(mem_41_2_R0_clk),
    .R0_data(mem_41_2_R0_data),
    .R0_en(mem_41_2_R0_en),
    .W0_addr(mem_41_2_W0_addr),
    .W0_clk(mem_41_2_W0_clk),
    .W0_data(mem_41_2_W0_data),
    .W0_en(mem_41_2_W0_en),
    .W0_mask(mem_41_2_W0_mask)
  );
  split_mem_0_ext mem_41_3 (
    .R0_addr(mem_41_3_R0_addr),
    .R0_clk(mem_41_3_R0_clk),
    .R0_data(mem_41_3_R0_data),
    .R0_en(mem_41_3_R0_en),
    .W0_addr(mem_41_3_W0_addr),
    .W0_clk(mem_41_3_W0_clk),
    .W0_data(mem_41_3_W0_data),
    .W0_en(mem_41_3_W0_en),
    .W0_mask(mem_41_3_W0_mask)
  );
  split_mem_0_ext mem_41_4 (
    .R0_addr(mem_41_4_R0_addr),
    .R0_clk(mem_41_4_R0_clk),
    .R0_data(mem_41_4_R0_data),
    .R0_en(mem_41_4_R0_en),
    .W0_addr(mem_41_4_W0_addr),
    .W0_clk(mem_41_4_W0_clk),
    .W0_data(mem_41_4_W0_data),
    .W0_en(mem_41_4_W0_en),
    .W0_mask(mem_41_4_W0_mask)
  );
  split_mem_0_ext mem_41_5 (
    .R0_addr(mem_41_5_R0_addr),
    .R0_clk(mem_41_5_R0_clk),
    .R0_data(mem_41_5_R0_data),
    .R0_en(mem_41_5_R0_en),
    .W0_addr(mem_41_5_W0_addr),
    .W0_clk(mem_41_5_W0_clk),
    .W0_data(mem_41_5_W0_data),
    .W0_en(mem_41_5_W0_en),
    .W0_mask(mem_41_5_W0_mask)
  );
  split_mem_0_ext mem_41_6 (
    .R0_addr(mem_41_6_R0_addr),
    .R0_clk(mem_41_6_R0_clk),
    .R0_data(mem_41_6_R0_data),
    .R0_en(mem_41_6_R0_en),
    .W0_addr(mem_41_6_W0_addr),
    .W0_clk(mem_41_6_W0_clk),
    .W0_data(mem_41_6_W0_data),
    .W0_en(mem_41_6_W0_en),
    .W0_mask(mem_41_6_W0_mask)
  );
  split_mem_0_ext mem_41_7 (
    .R0_addr(mem_41_7_R0_addr),
    .R0_clk(mem_41_7_R0_clk),
    .R0_data(mem_41_7_R0_data),
    .R0_en(mem_41_7_R0_en),
    .W0_addr(mem_41_7_W0_addr),
    .W0_clk(mem_41_7_W0_clk),
    .W0_data(mem_41_7_W0_data),
    .W0_en(mem_41_7_W0_en),
    .W0_mask(mem_41_7_W0_mask)
  );
  split_mem_0_ext mem_42_0 (
    .R0_addr(mem_42_0_R0_addr),
    .R0_clk(mem_42_0_R0_clk),
    .R0_data(mem_42_0_R0_data),
    .R0_en(mem_42_0_R0_en),
    .W0_addr(mem_42_0_W0_addr),
    .W0_clk(mem_42_0_W0_clk),
    .W0_data(mem_42_0_W0_data),
    .W0_en(mem_42_0_W0_en),
    .W0_mask(mem_42_0_W0_mask)
  );
  split_mem_0_ext mem_42_1 (
    .R0_addr(mem_42_1_R0_addr),
    .R0_clk(mem_42_1_R0_clk),
    .R0_data(mem_42_1_R0_data),
    .R0_en(mem_42_1_R0_en),
    .W0_addr(mem_42_1_W0_addr),
    .W0_clk(mem_42_1_W0_clk),
    .W0_data(mem_42_1_W0_data),
    .W0_en(mem_42_1_W0_en),
    .W0_mask(mem_42_1_W0_mask)
  );
  split_mem_0_ext mem_42_2 (
    .R0_addr(mem_42_2_R0_addr),
    .R0_clk(mem_42_2_R0_clk),
    .R0_data(mem_42_2_R0_data),
    .R0_en(mem_42_2_R0_en),
    .W0_addr(mem_42_2_W0_addr),
    .W0_clk(mem_42_2_W0_clk),
    .W0_data(mem_42_2_W0_data),
    .W0_en(mem_42_2_W0_en),
    .W0_mask(mem_42_2_W0_mask)
  );
  split_mem_0_ext mem_42_3 (
    .R0_addr(mem_42_3_R0_addr),
    .R0_clk(mem_42_3_R0_clk),
    .R0_data(mem_42_3_R0_data),
    .R0_en(mem_42_3_R0_en),
    .W0_addr(mem_42_3_W0_addr),
    .W0_clk(mem_42_3_W0_clk),
    .W0_data(mem_42_3_W0_data),
    .W0_en(mem_42_3_W0_en),
    .W0_mask(mem_42_3_W0_mask)
  );
  split_mem_0_ext mem_42_4 (
    .R0_addr(mem_42_4_R0_addr),
    .R0_clk(mem_42_4_R0_clk),
    .R0_data(mem_42_4_R0_data),
    .R0_en(mem_42_4_R0_en),
    .W0_addr(mem_42_4_W0_addr),
    .W0_clk(mem_42_4_W0_clk),
    .W0_data(mem_42_4_W0_data),
    .W0_en(mem_42_4_W0_en),
    .W0_mask(mem_42_4_W0_mask)
  );
  split_mem_0_ext mem_42_5 (
    .R0_addr(mem_42_5_R0_addr),
    .R0_clk(mem_42_5_R0_clk),
    .R0_data(mem_42_5_R0_data),
    .R0_en(mem_42_5_R0_en),
    .W0_addr(mem_42_5_W0_addr),
    .W0_clk(mem_42_5_W0_clk),
    .W0_data(mem_42_5_W0_data),
    .W0_en(mem_42_5_W0_en),
    .W0_mask(mem_42_5_W0_mask)
  );
  split_mem_0_ext mem_42_6 (
    .R0_addr(mem_42_6_R0_addr),
    .R0_clk(mem_42_6_R0_clk),
    .R0_data(mem_42_6_R0_data),
    .R0_en(mem_42_6_R0_en),
    .W0_addr(mem_42_6_W0_addr),
    .W0_clk(mem_42_6_W0_clk),
    .W0_data(mem_42_6_W0_data),
    .W0_en(mem_42_6_W0_en),
    .W0_mask(mem_42_6_W0_mask)
  );
  split_mem_0_ext mem_42_7 (
    .R0_addr(mem_42_7_R0_addr),
    .R0_clk(mem_42_7_R0_clk),
    .R0_data(mem_42_7_R0_data),
    .R0_en(mem_42_7_R0_en),
    .W0_addr(mem_42_7_W0_addr),
    .W0_clk(mem_42_7_W0_clk),
    .W0_data(mem_42_7_W0_data),
    .W0_en(mem_42_7_W0_en),
    .W0_mask(mem_42_7_W0_mask)
  );
  split_mem_0_ext mem_43_0 (
    .R0_addr(mem_43_0_R0_addr),
    .R0_clk(mem_43_0_R0_clk),
    .R0_data(mem_43_0_R0_data),
    .R0_en(mem_43_0_R0_en),
    .W0_addr(mem_43_0_W0_addr),
    .W0_clk(mem_43_0_W0_clk),
    .W0_data(mem_43_0_W0_data),
    .W0_en(mem_43_0_W0_en),
    .W0_mask(mem_43_0_W0_mask)
  );
  split_mem_0_ext mem_43_1 (
    .R0_addr(mem_43_1_R0_addr),
    .R0_clk(mem_43_1_R0_clk),
    .R0_data(mem_43_1_R0_data),
    .R0_en(mem_43_1_R0_en),
    .W0_addr(mem_43_1_W0_addr),
    .W0_clk(mem_43_1_W0_clk),
    .W0_data(mem_43_1_W0_data),
    .W0_en(mem_43_1_W0_en),
    .W0_mask(mem_43_1_W0_mask)
  );
  split_mem_0_ext mem_43_2 (
    .R0_addr(mem_43_2_R0_addr),
    .R0_clk(mem_43_2_R0_clk),
    .R0_data(mem_43_2_R0_data),
    .R0_en(mem_43_2_R0_en),
    .W0_addr(mem_43_2_W0_addr),
    .W0_clk(mem_43_2_W0_clk),
    .W0_data(mem_43_2_W0_data),
    .W0_en(mem_43_2_W0_en),
    .W0_mask(mem_43_2_W0_mask)
  );
  split_mem_0_ext mem_43_3 (
    .R0_addr(mem_43_3_R0_addr),
    .R0_clk(mem_43_3_R0_clk),
    .R0_data(mem_43_3_R0_data),
    .R0_en(mem_43_3_R0_en),
    .W0_addr(mem_43_3_W0_addr),
    .W0_clk(mem_43_3_W0_clk),
    .W0_data(mem_43_3_W0_data),
    .W0_en(mem_43_3_W0_en),
    .W0_mask(mem_43_3_W0_mask)
  );
  split_mem_0_ext mem_43_4 (
    .R0_addr(mem_43_4_R0_addr),
    .R0_clk(mem_43_4_R0_clk),
    .R0_data(mem_43_4_R0_data),
    .R0_en(mem_43_4_R0_en),
    .W0_addr(mem_43_4_W0_addr),
    .W0_clk(mem_43_4_W0_clk),
    .W0_data(mem_43_4_W0_data),
    .W0_en(mem_43_4_W0_en),
    .W0_mask(mem_43_4_W0_mask)
  );
  split_mem_0_ext mem_43_5 (
    .R0_addr(mem_43_5_R0_addr),
    .R0_clk(mem_43_5_R0_clk),
    .R0_data(mem_43_5_R0_data),
    .R0_en(mem_43_5_R0_en),
    .W0_addr(mem_43_5_W0_addr),
    .W0_clk(mem_43_5_W0_clk),
    .W0_data(mem_43_5_W0_data),
    .W0_en(mem_43_5_W0_en),
    .W0_mask(mem_43_5_W0_mask)
  );
  split_mem_0_ext mem_43_6 (
    .R0_addr(mem_43_6_R0_addr),
    .R0_clk(mem_43_6_R0_clk),
    .R0_data(mem_43_6_R0_data),
    .R0_en(mem_43_6_R0_en),
    .W0_addr(mem_43_6_W0_addr),
    .W0_clk(mem_43_6_W0_clk),
    .W0_data(mem_43_6_W0_data),
    .W0_en(mem_43_6_W0_en),
    .W0_mask(mem_43_6_W0_mask)
  );
  split_mem_0_ext mem_43_7 (
    .R0_addr(mem_43_7_R0_addr),
    .R0_clk(mem_43_7_R0_clk),
    .R0_data(mem_43_7_R0_data),
    .R0_en(mem_43_7_R0_en),
    .W0_addr(mem_43_7_W0_addr),
    .W0_clk(mem_43_7_W0_clk),
    .W0_data(mem_43_7_W0_data),
    .W0_en(mem_43_7_W0_en),
    .W0_mask(mem_43_7_W0_mask)
  );
  split_mem_0_ext mem_44_0 (
    .R0_addr(mem_44_0_R0_addr),
    .R0_clk(mem_44_0_R0_clk),
    .R0_data(mem_44_0_R0_data),
    .R0_en(mem_44_0_R0_en),
    .W0_addr(mem_44_0_W0_addr),
    .W0_clk(mem_44_0_W0_clk),
    .W0_data(mem_44_0_W0_data),
    .W0_en(mem_44_0_W0_en),
    .W0_mask(mem_44_0_W0_mask)
  );
  split_mem_0_ext mem_44_1 (
    .R0_addr(mem_44_1_R0_addr),
    .R0_clk(mem_44_1_R0_clk),
    .R0_data(mem_44_1_R0_data),
    .R0_en(mem_44_1_R0_en),
    .W0_addr(mem_44_1_W0_addr),
    .W0_clk(mem_44_1_W0_clk),
    .W0_data(mem_44_1_W0_data),
    .W0_en(mem_44_1_W0_en),
    .W0_mask(mem_44_1_W0_mask)
  );
  split_mem_0_ext mem_44_2 (
    .R0_addr(mem_44_2_R0_addr),
    .R0_clk(mem_44_2_R0_clk),
    .R0_data(mem_44_2_R0_data),
    .R0_en(mem_44_2_R0_en),
    .W0_addr(mem_44_2_W0_addr),
    .W0_clk(mem_44_2_W0_clk),
    .W0_data(mem_44_2_W0_data),
    .W0_en(mem_44_2_W0_en),
    .W0_mask(mem_44_2_W0_mask)
  );
  split_mem_0_ext mem_44_3 (
    .R0_addr(mem_44_3_R0_addr),
    .R0_clk(mem_44_3_R0_clk),
    .R0_data(mem_44_3_R0_data),
    .R0_en(mem_44_3_R0_en),
    .W0_addr(mem_44_3_W0_addr),
    .W0_clk(mem_44_3_W0_clk),
    .W0_data(mem_44_3_W0_data),
    .W0_en(mem_44_3_W0_en),
    .W0_mask(mem_44_3_W0_mask)
  );
  split_mem_0_ext mem_44_4 (
    .R0_addr(mem_44_4_R0_addr),
    .R0_clk(mem_44_4_R0_clk),
    .R0_data(mem_44_4_R0_data),
    .R0_en(mem_44_4_R0_en),
    .W0_addr(mem_44_4_W0_addr),
    .W0_clk(mem_44_4_W0_clk),
    .W0_data(mem_44_4_W0_data),
    .W0_en(mem_44_4_W0_en),
    .W0_mask(mem_44_4_W0_mask)
  );
  split_mem_0_ext mem_44_5 (
    .R0_addr(mem_44_5_R0_addr),
    .R0_clk(mem_44_5_R0_clk),
    .R0_data(mem_44_5_R0_data),
    .R0_en(mem_44_5_R0_en),
    .W0_addr(mem_44_5_W0_addr),
    .W0_clk(mem_44_5_W0_clk),
    .W0_data(mem_44_5_W0_data),
    .W0_en(mem_44_5_W0_en),
    .W0_mask(mem_44_5_W0_mask)
  );
  split_mem_0_ext mem_44_6 (
    .R0_addr(mem_44_6_R0_addr),
    .R0_clk(mem_44_6_R0_clk),
    .R0_data(mem_44_6_R0_data),
    .R0_en(mem_44_6_R0_en),
    .W0_addr(mem_44_6_W0_addr),
    .W0_clk(mem_44_6_W0_clk),
    .W0_data(mem_44_6_W0_data),
    .W0_en(mem_44_6_W0_en),
    .W0_mask(mem_44_6_W0_mask)
  );
  split_mem_0_ext mem_44_7 (
    .R0_addr(mem_44_7_R0_addr),
    .R0_clk(mem_44_7_R0_clk),
    .R0_data(mem_44_7_R0_data),
    .R0_en(mem_44_7_R0_en),
    .W0_addr(mem_44_7_W0_addr),
    .W0_clk(mem_44_7_W0_clk),
    .W0_data(mem_44_7_W0_data),
    .W0_en(mem_44_7_W0_en),
    .W0_mask(mem_44_7_W0_mask)
  );
  split_mem_0_ext mem_45_0 (
    .R0_addr(mem_45_0_R0_addr),
    .R0_clk(mem_45_0_R0_clk),
    .R0_data(mem_45_0_R0_data),
    .R0_en(mem_45_0_R0_en),
    .W0_addr(mem_45_0_W0_addr),
    .W0_clk(mem_45_0_W0_clk),
    .W0_data(mem_45_0_W0_data),
    .W0_en(mem_45_0_W0_en),
    .W0_mask(mem_45_0_W0_mask)
  );
  split_mem_0_ext mem_45_1 (
    .R0_addr(mem_45_1_R0_addr),
    .R0_clk(mem_45_1_R0_clk),
    .R0_data(mem_45_1_R0_data),
    .R0_en(mem_45_1_R0_en),
    .W0_addr(mem_45_1_W0_addr),
    .W0_clk(mem_45_1_W0_clk),
    .W0_data(mem_45_1_W0_data),
    .W0_en(mem_45_1_W0_en),
    .W0_mask(mem_45_1_W0_mask)
  );
  split_mem_0_ext mem_45_2 (
    .R0_addr(mem_45_2_R0_addr),
    .R0_clk(mem_45_2_R0_clk),
    .R0_data(mem_45_2_R0_data),
    .R0_en(mem_45_2_R0_en),
    .W0_addr(mem_45_2_W0_addr),
    .W0_clk(mem_45_2_W0_clk),
    .W0_data(mem_45_2_W0_data),
    .W0_en(mem_45_2_W0_en),
    .W0_mask(mem_45_2_W0_mask)
  );
  split_mem_0_ext mem_45_3 (
    .R0_addr(mem_45_3_R0_addr),
    .R0_clk(mem_45_3_R0_clk),
    .R0_data(mem_45_3_R0_data),
    .R0_en(mem_45_3_R0_en),
    .W0_addr(mem_45_3_W0_addr),
    .W0_clk(mem_45_3_W0_clk),
    .W0_data(mem_45_3_W0_data),
    .W0_en(mem_45_3_W0_en),
    .W0_mask(mem_45_3_W0_mask)
  );
  split_mem_0_ext mem_45_4 (
    .R0_addr(mem_45_4_R0_addr),
    .R0_clk(mem_45_4_R0_clk),
    .R0_data(mem_45_4_R0_data),
    .R0_en(mem_45_4_R0_en),
    .W0_addr(mem_45_4_W0_addr),
    .W0_clk(mem_45_4_W0_clk),
    .W0_data(mem_45_4_W0_data),
    .W0_en(mem_45_4_W0_en),
    .W0_mask(mem_45_4_W0_mask)
  );
  split_mem_0_ext mem_45_5 (
    .R0_addr(mem_45_5_R0_addr),
    .R0_clk(mem_45_5_R0_clk),
    .R0_data(mem_45_5_R0_data),
    .R0_en(mem_45_5_R0_en),
    .W0_addr(mem_45_5_W0_addr),
    .W0_clk(mem_45_5_W0_clk),
    .W0_data(mem_45_5_W0_data),
    .W0_en(mem_45_5_W0_en),
    .W0_mask(mem_45_5_W0_mask)
  );
  split_mem_0_ext mem_45_6 (
    .R0_addr(mem_45_6_R0_addr),
    .R0_clk(mem_45_6_R0_clk),
    .R0_data(mem_45_6_R0_data),
    .R0_en(mem_45_6_R0_en),
    .W0_addr(mem_45_6_W0_addr),
    .W0_clk(mem_45_6_W0_clk),
    .W0_data(mem_45_6_W0_data),
    .W0_en(mem_45_6_W0_en),
    .W0_mask(mem_45_6_W0_mask)
  );
  split_mem_0_ext mem_45_7 (
    .R0_addr(mem_45_7_R0_addr),
    .R0_clk(mem_45_7_R0_clk),
    .R0_data(mem_45_7_R0_data),
    .R0_en(mem_45_7_R0_en),
    .W0_addr(mem_45_7_W0_addr),
    .W0_clk(mem_45_7_W0_clk),
    .W0_data(mem_45_7_W0_data),
    .W0_en(mem_45_7_W0_en),
    .W0_mask(mem_45_7_W0_mask)
  );
  split_mem_0_ext mem_46_0 (
    .R0_addr(mem_46_0_R0_addr),
    .R0_clk(mem_46_0_R0_clk),
    .R0_data(mem_46_0_R0_data),
    .R0_en(mem_46_0_R0_en),
    .W0_addr(mem_46_0_W0_addr),
    .W0_clk(mem_46_0_W0_clk),
    .W0_data(mem_46_0_W0_data),
    .W0_en(mem_46_0_W0_en),
    .W0_mask(mem_46_0_W0_mask)
  );
  split_mem_0_ext mem_46_1 (
    .R0_addr(mem_46_1_R0_addr),
    .R0_clk(mem_46_1_R0_clk),
    .R0_data(mem_46_1_R0_data),
    .R0_en(mem_46_1_R0_en),
    .W0_addr(mem_46_1_W0_addr),
    .W0_clk(mem_46_1_W0_clk),
    .W0_data(mem_46_1_W0_data),
    .W0_en(mem_46_1_W0_en),
    .W0_mask(mem_46_1_W0_mask)
  );
  split_mem_0_ext mem_46_2 (
    .R0_addr(mem_46_2_R0_addr),
    .R0_clk(mem_46_2_R0_clk),
    .R0_data(mem_46_2_R0_data),
    .R0_en(mem_46_2_R0_en),
    .W0_addr(mem_46_2_W0_addr),
    .W0_clk(mem_46_2_W0_clk),
    .W0_data(mem_46_2_W0_data),
    .W0_en(mem_46_2_W0_en),
    .W0_mask(mem_46_2_W0_mask)
  );
  split_mem_0_ext mem_46_3 (
    .R0_addr(mem_46_3_R0_addr),
    .R0_clk(mem_46_3_R0_clk),
    .R0_data(mem_46_3_R0_data),
    .R0_en(mem_46_3_R0_en),
    .W0_addr(mem_46_3_W0_addr),
    .W0_clk(mem_46_3_W0_clk),
    .W0_data(mem_46_3_W0_data),
    .W0_en(mem_46_3_W0_en),
    .W0_mask(mem_46_3_W0_mask)
  );
  split_mem_0_ext mem_46_4 (
    .R0_addr(mem_46_4_R0_addr),
    .R0_clk(mem_46_4_R0_clk),
    .R0_data(mem_46_4_R0_data),
    .R0_en(mem_46_4_R0_en),
    .W0_addr(mem_46_4_W0_addr),
    .W0_clk(mem_46_4_W0_clk),
    .W0_data(mem_46_4_W0_data),
    .W0_en(mem_46_4_W0_en),
    .W0_mask(mem_46_4_W0_mask)
  );
  split_mem_0_ext mem_46_5 (
    .R0_addr(mem_46_5_R0_addr),
    .R0_clk(mem_46_5_R0_clk),
    .R0_data(mem_46_5_R0_data),
    .R0_en(mem_46_5_R0_en),
    .W0_addr(mem_46_5_W0_addr),
    .W0_clk(mem_46_5_W0_clk),
    .W0_data(mem_46_5_W0_data),
    .W0_en(mem_46_5_W0_en),
    .W0_mask(mem_46_5_W0_mask)
  );
  split_mem_0_ext mem_46_6 (
    .R0_addr(mem_46_6_R0_addr),
    .R0_clk(mem_46_6_R0_clk),
    .R0_data(mem_46_6_R0_data),
    .R0_en(mem_46_6_R0_en),
    .W0_addr(mem_46_6_W0_addr),
    .W0_clk(mem_46_6_W0_clk),
    .W0_data(mem_46_6_W0_data),
    .W0_en(mem_46_6_W0_en),
    .W0_mask(mem_46_6_W0_mask)
  );
  split_mem_0_ext mem_46_7 (
    .R0_addr(mem_46_7_R0_addr),
    .R0_clk(mem_46_7_R0_clk),
    .R0_data(mem_46_7_R0_data),
    .R0_en(mem_46_7_R0_en),
    .W0_addr(mem_46_7_W0_addr),
    .W0_clk(mem_46_7_W0_clk),
    .W0_data(mem_46_7_W0_data),
    .W0_en(mem_46_7_W0_en),
    .W0_mask(mem_46_7_W0_mask)
  );
  split_mem_0_ext mem_47_0 (
    .R0_addr(mem_47_0_R0_addr),
    .R0_clk(mem_47_0_R0_clk),
    .R0_data(mem_47_0_R0_data),
    .R0_en(mem_47_0_R0_en),
    .W0_addr(mem_47_0_W0_addr),
    .W0_clk(mem_47_0_W0_clk),
    .W0_data(mem_47_0_W0_data),
    .W0_en(mem_47_0_W0_en),
    .W0_mask(mem_47_0_W0_mask)
  );
  split_mem_0_ext mem_47_1 (
    .R0_addr(mem_47_1_R0_addr),
    .R0_clk(mem_47_1_R0_clk),
    .R0_data(mem_47_1_R0_data),
    .R0_en(mem_47_1_R0_en),
    .W0_addr(mem_47_1_W0_addr),
    .W0_clk(mem_47_1_W0_clk),
    .W0_data(mem_47_1_W0_data),
    .W0_en(mem_47_1_W0_en),
    .W0_mask(mem_47_1_W0_mask)
  );
  split_mem_0_ext mem_47_2 (
    .R0_addr(mem_47_2_R0_addr),
    .R0_clk(mem_47_2_R0_clk),
    .R0_data(mem_47_2_R0_data),
    .R0_en(mem_47_2_R0_en),
    .W0_addr(mem_47_2_W0_addr),
    .W0_clk(mem_47_2_W0_clk),
    .W0_data(mem_47_2_W0_data),
    .W0_en(mem_47_2_W0_en),
    .W0_mask(mem_47_2_W0_mask)
  );
  split_mem_0_ext mem_47_3 (
    .R0_addr(mem_47_3_R0_addr),
    .R0_clk(mem_47_3_R0_clk),
    .R0_data(mem_47_3_R0_data),
    .R0_en(mem_47_3_R0_en),
    .W0_addr(mem_47_3_W0_addr),
    .W0_clk(mem_47_3_W0_clk),
    .W0_data(mem_47_3_W0_data),
    .W0_en(mem_47_3_W0_en),
    .W0_mask(mem_47_3_W0_mask)
  );
  split_mem_0_ext mem_47_4 (
    .R0_addr(mem_47_4_R0_addr),
    .R0_clk(mem_47_4_R0_clk),
    .R0_data(mem_47_4_R0_data),
    .R0_en(mem_47_4_R0_en),
    .W0_addr(mem_47_4_W0_addr),
    .W0_clk(mem_47_4_W0_clk),
    .W0_data(mem_47_4_W0_data),
    .W0_en(mem_47_4_W0_en),
    .W0_mask(mem_47_4_W0_mask)
  );
  split_mem_0_ext mem_47_5 (
    .R0_addr(mem_47_5_R0_addr),
    .R0_clk(mem_47_5_R0_clk),
    .R0_data(mem_47_5_R0_data),
    .R0_en(mem_47_5_R0_en),
    .W0_addr(mem_47_5_W0_addr),
    .W0_clk(mem_47_5_W0_clk),
    .W0_data(mem_47_5_W0_data),
    .W0_en(mem_47_5_W0_en),
    .W0_mask(mem_47_5_W0_mask)
  );
  split_mem_0_ext mem_47_6 (
    .R0_addr(mem_47_6_R0_addr),
    .R0_clk(mem_47_6_R0_clk),
    .R0_data(mem_47_6_R0_data),
    .R0_en(mem_47_6_R0_en),
    .W0_addr(mem_47_6_W0_addr),
    .W0_clk(mem_47_6_W0_clk),
    .W0_data(mem_47_6_W0_data),
    .W0_en(mem_47_6_W0_en),
    .W0_mask(mem_47_6_W0_mask)
  );
  split_mem_0_ext mem_47_7 (
    .R0_addr(mem_47_7_R0_addr),
    .R0_clk(mem_47_7_R0_clk),
    .R0_data(mem_47_7_R0_data),
    .R0_en(mem_47_7_R0_en),
    .W0_addr(mem_47_7_W0_addr),
    .W0_clk(mem_47_7_W0_clk),
    .W0_data(mem_47_7_W0_data),
    .W0_en(mem_47_7_W0_en),
    .W0_mask(mem_47_7_W0_mask)
  );
  split_mem_0_ext mem_48_0 (
    .R0_addr(mem_48_0_R0_addr),
    .R0_clk(mem_48_0_R0_clk),
    .R0_data(mem_48_0_R0_data),
    .R0_en(mem_48_0_R0_en),
    .W0_addr(mem_48_0_W0_addr),
    .W0_clk(mem_48_0_W0_clk),
    .W0_data(mem_48_0_W0_data),
    .W0_en(mem_48_0_W0_en),
    .W0_mask(mem_48_0_W0_mask)
  );
  split_mem_0_ext mem_48_1 (
    .R0_addr(mem_48_1_R0_addr),
    .R0_clk(mem_48_1_R0_clk),
    .R0_data(mem_48_1_R0_data),
    .R0_en(mem_48_1_R0_en),
    .W0_addr(mem_48_1_W0_addr),
    .W0_clk(mem_48_1_W0_clk),
    .W0_data(mem_48_1_W0_data),
    .W0_en(mem_48_1_W0_en),
    .W0_mask(mem_48_1_W0_mask)
  );
  split_mem_0_ext mem_48_2 (
    .R0_addr(mem_48_2_R0_addr),
    .R0_clk(mem_48_2_R0_clk),
    .R0_data(mem_48_2_R0_data),
    .R0_en(mem_48_2_R0_en),
    .W0_addr(mem_48_2_W0_addr),
    .W0_clk(mem_48_2_W0_clk),
    .W0_data(mem_48_2_W0_data),
    .W0_en(mem_48_2_W0_en),
    .W0_mask(mem_48_2_W0_mask)
  );
  split_mem_0_ext mem_48_3 (
    .R0_addr(mem_48_3_R0_addr),
    .R0_clk(mem_48_3_R0_clk),
    .R0_data(mem_48_3_R0_data),
    .R0_en(mem_48_3_R0_en),
    .W0_addr(mem_48_3_W0_addr),
    .W0_clk(mem_48_3_W0_clk),
    .W0_data(mem_48_3_W0_data),
    .W0_en(mem_48_3_W0_en),
    .W0_mask(mem_48_3_W0_mask)
  );
  split_mem_0_ext mem_48_4 (
    .R0_addr(mem_48_4_R0_addr),
    .R0_clk(mem_48_4_R0_clk),
    .R0_data(mem_48_4_R0_data),
    .R0_en(mem_48_4_R0_en),
    .W0_addr(mem_48_4_W0_addr),
    .W0_clk(mem_48_4_W0_clk),
    .W0_data(mem_48_4_W0_data),
    .W0_en(mem_48_4_W0_en),
    .W0_mask(mem_48_4_W0_mask)
  );
  split_mem_0_ext mem_48_5 (
    .R0_addr(mem_48_5_R0_addr),
    .R0_clk(mem_48_5_R0_clk),
    .R0_data(mem_48_5_R0_data),
    .R0_en(mem_48_5_R0_en),
    .W0_addr(mem_48_5_W0_addr),
    .W0_clk(mem_48_5_W0_clk),
    .W0_data(mem_48_5_W0_data),
    .W0_en(mem_48_5_W0_en),
    .W0_mask(mem_48_5_W0_mask)
  );
  split_mem_0_ext mem_48_6 (
    .R0_addr(mem_48_6_R0_addr),
    .R0_clk(mem_48_6_R0_clk),
    .R0_data(mem_48_6_R0_data),
    .R0_en(mem_48_6_R0_en),
    .W0_addr(mem_48_6_W0_addr),
    .W0_clk(mem_48_6_W0_clk),
    .W0_data(mem_48_6_W0_data),
    .W0_en(mem_48_6_W0_en),
    .W0_mask(mem_48_6_W0_mask)
  );
  split_mem_0_ext mem_48_7 (
    .R0_addr(mem_48_7_R0_addr),
    .R0_clk(mem_48_7_R0_clk),
    .R0_data(mem_48_7_R0_data),
    .R0_en(mem_48_7_R0_en),
    .W0_addr(mem_48_7_W0_addr),
    .W0_clk(mem_48_7_W0_clk),
    .W0_data(mem_48_7_W0_data),
    .W0_en(mem_48_7_W0_en),
    .W0_mask(mem_48_7_W0_mask)
  );
  split_mem_0_ext mem_49_0 (
    .R0_addr(mem_49_0_R0_addr),
    .R0_clk(mem_49_0_R0_clk),
    .R0_data(mem_49_0_R0_data),
    .R0_en(mem_49_0_R0_en),
    .W0_addr(mem_49_0_W0_addr),
    .W0_clk(mem_49_0_W0_clk),
    .W0_data(mem_49_0_W0_data),
    .W0_en(mem_49_0_W0_en),
    .W0_mask(mem_49_0_W0_mask)
  );
  split_mem_0_ext mem_49_1 (
    .R0_addr(mem_49_1_R0_addr),
    .R0_clk(mem_49_1_R0_clk),
    .R0_data(mem_49_1_R0_data),
    .R0_en(mem_49_1_R0_en),
    .W0_addr(mem_49_1_W0_addr),
    .W0_clk(mem_49_1_W0_clk),
    .W0_data(mem_49_1_W0_data),
    .W0_en(mem_49_1_W0_en),
    .W0_mask(mem_49_1_W0_mask)
  );
  split_mem_0_ext mem_49_2 (
    .R0_addr(mem_49_2_R0_addr),
    .R0_clk(mem_49_2_R0_clk),
    .R0_data(mem_49_2_R0_data),
    .R0_en(mem_49_2_R0_en),
    .W0_addr(mem_49_2_W0_addr),
    .W0_clk(mem_49_2_W0_clk),
    .W0_data(mem_49_2_W0_data),
    .W0_en(mem_49_2_W0_en),
    .W0_mask(mem_49_2_W0_mask)
  );
  split_mem_0_ext mem_49_3 (
    .R0_addr(mem_49_3_R0_addr),
    .R0_clk(mem_49_3_R0_clk),
    .R0_data(mem_49_3_R0_data),
    .R0_en(mem_49_3_R0_en),
    .W0_addr(mem_49_3_W0_addr),
    .W0_clk(mem_49_3_W0_clk),
    .W0_data(mem_49_3_W0_data),
    .W0_en(mem_49_3_W0_en),
    .W0_mask(mem_49_3_W0_mask)
  );
  split_mem_0_ext mem_49_4 (
    .R0_addr(mem_49_4_R0_addr),
    .R0_clk(mem_49_4_R0_clk),
    .R0_data(mem_49_4_R0_data),
    .R0_en(mem_49_4_R0_en),
    .W0_addr(mem_49_4_W0_addr),
    .W0_clk(mem_49_4_W0_clk),
    .W0_data(mem_49_4_W0_data),
    .W0_en(mem_49_4_W0_en),
    .W0_mask(mem_49_4_W0_mask)
  );
  split_mem_0_ext mem_49_5 (
    .R0_addr(mem_49_5_R0_addr),
    .R0_clk(mem_49_5_R0_clk),
    .R0_data(mem_49_5_R0_data),
    .R0_en(mem_49_5_R0_en),
    .W0_addr(mem_49_5_W0_addr),
    .W0_clk(mem_49_5_W0_clk),
    .W0_data(mem_49_5_W0_data),
    .W0_en(mem_49_5_W0_en),
    .W0_mask(mem_49_5_W0_mask)
  );
  split_mem_0_ext mem_49_6 (
    .R0_addr(mem_49_6_R0_addr),
    .R0_clk(mem_49_6_R0_clk),
    .R0_data(mem_49_6_R0_data),
    .R0_en(mem_49_6_R0_en),
    .W0_addr(mem_49_6_W0_addr),
    .W0_clk(mem_49_6_W0_clk),
    .W0_data(mem_49_6_W0_data),
    .W0_en(mem_49_6_W0_en),
    .W0_mask(mem_49_6_W0_mask)
  );
  split_mem_0_ext mem_49_7 (
    .R0_addr(mem_49_7_R0_addr),
    .R0_clk(mem_49_7_R0_clk),
    .R0_data(mem_49_7_R0_data),
    .R0_en(mem_49_7_R0_en),
    .W0_addr(mem_49_7_W0_addr),
    .W0_clk(mem_49_7_W0_clk),
    .W0_data(mem_49_7_W0_data),
    .W0_en(mem_49_7_W0_en),
    .W0_mask(mem_49_7_W0_mask)
  );
  split_mem_0_ext mem_50_0 (
    .R0_addr(mem_50_0_R0_addr),
    .R0_clk(mem_50_0_R0_clk),
    .R0_data(mem_50_0_R0_data),
    .R0_en(mem_50_0_R0_en),
    .W0_addr(mem_50_0_W0_addr),
    .W0_clk(mem_50_0_W0_clk),
    .W0_data(mem_50_0_W0_data),
    .W0_en(mem_50_0_W0_en),
    .W0_mask(mem_50_0_W0_mask)
  );
  split_mem_0_ext mem_50_1 (
    .R0_addr(mem_50_1_R0_addr),
    .R0_clk(mem_50_1_R0_clk),
    .R0_data(mem_50_1_R0_data),
    .R0_en(mem_50_1_R0_en),
    .W0_addr(mem_50_1_W0_addr),
    .W0_clk(mem_50_1_W0_clk),
    .W0_data(mem_50_1_W0_data),
    .W0_en(mem_50_1_W0_en),
    .W0_mask(mem_50_1_W0_mask)
  );
  split_mem_0_ext mem_50_2 (
    .R0_addr(mem_50_2_R0_addr),
    .R0_clk(mem_50_2_R0_clk),
    .R0_data(mem_50_2_R0_data),
    .R0_en(mem_50_2_R0_en),
    .W0_addr(mem_50_2_W0_addr),
    .W0_clk(mem_50_2_W0_clk),
    .W0_data(mem_50_2_W0_data),
    .W0_en(mem_50_2_W0_en),
    .W0_mask(mem_50_2_W0_mask)
  );
  split_mem_0_ext mem_50_3 (
    .R0_addr(mem_50_3_R0_addr),
    .R0_clk(mem_50_3_R0_clk),
    .R0_data(mem_50_3_R0_data),
    .R0_en(mem_50_3_R0_en),
    .W0_addr(mem_50_3_W0_addr),
    .W0_clk(mem_50_3_W0_clk),
    .W0_data(mem_50_3_W0_data),
    .W0_en(mem_50_3_W0_en),
    .W0_mask(mem_50_3_W0_mask)
  );
  split_mem_0_ext mem_50_4 (
    .R0_addr(mem_50_4_R0_addr),
    .R0_clk(mem_50_4_R0_clk),
    .R0_data(mem_50_4_R0_data),
    .R0_en(mem_50_4_R0_en),
    .W0_addr(mem_50_4_W0_addr),
    .W0_clk(mem_50_4_W0_clk),
    .W0_data(mem_50_4_W0_data),
    .W0_en(mem_50_4_W0_en),
    .W0_mask(mem_50_4_W0_mask)
  );
  split_mem_0_ext mem_50_5 (
    .R0_addr(mem_50_5_R0_addr),
    .R0_clk(mem_50_5_R0_clk),
    .R0_data(mem_50_5_R0_data),
    .R0_en(mem_50_5_R0_en),
    .W0_addr(mem_50_5_W0_addr),
    .W0_clk(mem_50_5_W0_clk),
    .W0_data(mem_50_5_W0_data),
    .W0_en(mem_50_5_W0_en),
    .W0_mask(mem_50_5_W0_mask)
  );
  split_mem_0_ext mem_50_6 (
    .R0_addr(mem_50_6_R0_addr),
    .R0_clk(mem_50_6_R0_clk),
    .R0_data(mem_50_6_R0_data),
    .R0_en(mem_50_6_R0_en),
    .W0_addr(mem_50_6_W0_addr),
    .W0_clk(mem_50_6_W0_clk),
    .W0_data(mem_50_6_W0_data),
    .W0_en(mem_50_6_W0_en),
    .W0_mask(mem_50_6_W0_mask)
  );
  split_mem_0_ext mem_50_7 (
    .R0_addr(mem_50_7_R0_addr),
    .R0_clk(mem_50_7_R0_clk),
    .R0_data(mem_50_7_R0_data),
    .R0_en(mem_50_7_R0_en),
    .W0_addr(mem_50_7_W0_addr),
    .W0_clk(mem_50_7_W0_clk),
    .W0_data(mem_50_7_W0_data),
    .W0_en(mem_50_7_W0_en),
    .W0_mask(mem_50_7_W0_mask)
  );
  split_mem_0_ext mem_51_0 (
    .R0_addr(mem_51_0_R0_addr),
    .R0_clk(mem_51_0_R0_clk),
    .R0_data(mem_51_0_R0_data),
    .R0_en(mem_51_0_R0_en),
    .W0_addr(mem_51_0_W0_addr),
    .W0_clk(mem_51_0_W0_clk),
    .W0_data(mem_51_0_W0_data),
    .W0_en(mem_51_0_W0_en),
    .W0_mask(mem_51_0_W0_mask)
  );
  split_mem_0_ext mem_51_1 (
    .R0_addr(mem_51_1_R0_addr),
    .R0_clk(mem_51_1_R0_clk),
    .R0_data(mem_51_1_R0_data),
    .R0_en(mem_51_1_R0_en),
    .W0_addr(mem_51_1_W0_addr),
    .W0_clk(mem_51_1_W0_clk),
    .W0_data(mem_51_1_W0_data),
    .W0_en(mem_51_1_W0_en),
    .W0_mask(mem_51_1_W0_mask)
  );
  split_mem_0_ext mem_51_2 (
    .R0_addr(mem_51_2_R0_addr),
    .R0_clk(mem_51_2_R0_clk),
    .R0_data(mem_51_2_R0_data),
    .R0_en(mem_51_2_R0_en),
    .W0_addr(mem_51_2_W0_addr),
    .W0_clk(mem_51_2_W0_clk),
    .W0_data(mem_51_2_W0_data),
    .W0_en(mem_51_2_W0_en),
    .W0_mask(mem_51_2_W0_mask)
  );
  split_mem_0_ext mem_51_3 (
    .R0_addr(mem_51_3_R0_addr),
    .R0_clk(mem_51_3_R0_clk),
    .R0_data(mem_51_3_R0_data),
    .R0_en(mem_51_3_R0_en),
    .W0_addr(mem_51_3_W0_addr),
    .W0_clk(mem_51_3_W0_clk),
    .W0_data(mem_51_3_W0_data),
    .W0_en(mem_51_3_W0_en),
    .W0_mask(mem_51_3_W0_mask)
  );
  split_mem_0_ext mem_51_4 (
    .R0_addr(mem_51_4_R0_addr),
    .R0_clk(mem_51_4_R0_clk),
    .R0_data(mem_51_4_R0_data),
    .R0_en(mem_51_4_R0_en),
    .W0_addr(mem_51_4_W0_addr),
    .W0_clk(mem_51_4_W0_clk),
    .W0_data(mem_51_4_W0_data),
    .W0_en(mem_51_4_W0_en),
    .W0_mask(mem_51_4_W0_mask)
  );
  split_mem_0_ext mem_51_5 (
    .R0_addr(mem_51_5_R0_addr),
    .R0_clk(mem_51_5_R0_clk),
    .R0_data(mem_51_5_R0_data),
    .R0_en(mem_51_5_R0_en),
    .W0_addr(mem_51_5_W0_addr),
    .W0_clk(mem_51_5_W0_clk),
    .W0_data(mem_51_5_W0_data),
    .W0_en(mem_51_5_W0_en),
    .W0_mask(mem_51_5_W0_mask)
  );
  split_mem_0_ext mem_51_6 (
    .R0_addr(mem_51_6_R0_addr),
    .R0_clk(mem_51_6_R0_clk),
    .R0_data(mem_51_6_R0_data),
    .R0_en(mem_51_6_R0_en),
    .W0_addr(mem_51_6_W0_addr),
    .W0_clk(mem_51_6_W0_clk),
    .W0_data(mem_51_6_W0_data),
    .W0_en(mem_51_6_W0_en),
    .W0_mask(mem_51_6_W0_mask)
  );
  split_mem_0_ext mem_51_7 (
    .R0_addr(mem_51_7_R0_addr),
    .R0_clk(mem_51_7_R0_clk),
    .R0_data(mem_51_7_R0_data),
    .R0_en(mem_51_7_R0_en),
    .W0_addr(mem_51_7_W0_addr),
    .W0_clk(mem_51_7_W0_clk),
    .W0_data(mem_51_7_W0_data),
    .W0_en(mem_51_7_W0_en),
    .W0_mask(mem_51_7_W0_mask)
  );
  split_mem_0_ext mem_52_0 (
    .R0_addr(mem_52_0_R0_addr),
    .R0_clk(mem_52_0_R0_clk),
    .R0_data(mem_52_0_R0_data),
    .R0_en(mem_52_0_R0_en),
    .W0_addr(mem_52_0_W0_addr),
    .W0_clk(mem_52_0_W0_clk),
    .W0_data(mem_52_0_W0_data),
    .W0_en(mem_52_0_W0_en),
    .W0_mask(mem_52_0_W0_mask)
  );
  split_mem_0_ext mem_52_1 (
    .R0_addr(mem_52_1_R0_addr),
    .R0_clk(mem_52_1_R0_clk),
    .R0_data(mem_52_1_R0_data),
    .R0_en(mem_52_1_R0_en),
    .W0_addr(mem_52_1_W0_addr),
    .W0_clk(mem_52_1_W0_clk),
    .W0_data(mem_52_1_W0_data),
    .W0_en(mem_52_1_W0_en),
    .W0_mask(mem_52_1_W0_mask)
  );
  split_mem_0_ext mem_52_2 (
    .R0_addr(mem_52_2_R0_addr),
    .R0_clk(mem_52_2_R0_clk),
    .R0_data(mem_52_2_R0_data),
    .R0_en(mem_52_2_R0_en),
    .W0_addr(mem_52_2_W0_addr),
    .W0_clk(mem_52_2_W0_clk),
    .W0_data(mem_52_2_W0_data),
    .W0_en(mem_52_2_W0_en),
    .W0_mask(mem_52_2_W0_mask)
  );
  split_mem_0_ext mem_52_3 (
    .R0_addr(mem_52_3_R0_addr),
    .R0_clk(mem_52_3_R0_clk),
    .R0_data(mem_52_3_R0_data),
    .R0_en(mem_52_3_R0_en),
    .W0_addr(mem_52_3_W0_addr),
    .W0_clk(mem_52_3_W0_clk),
    .W0_data(mem_52_3_W0_data),
    .W0_en(mem_52_3_W0_en),
    .W0_mask(mem_52_3_W0_mask)
  );
  split_mem_0_ext mem_52_4 (
    .R0_addr(mem_52_4_R0_addr),
    .R0_clk(mem_52_4_R0_clk),
    .R0_data(mem_52_4_R0_data),
    .R0_en(mem_52_4_R0_en),
    .W0_addr(mem_52_4_W0_addr),
    .W0_clk(mem_52_4_W0_clk),
    .W0_data(mem_52_4_W0_data),
    .W0_en(mem_52_4_W0_en),
    .W0_mask(mem_52_4_W0_mask)
  );
  split_mem_0_ext mem_52_5 (
    .R0_addr(mem_52_5_R0_addr),
    .R0_clk(mem_52_5_R0_clk),
    .R0_data(mem_52_5_R0_data),
    .R0_en(mem_52_5_R0_en),
    .W0_addr(mem_52_5_W0_addr),
    .W0_clk(mem_52_5_W0_clk),
    .W0_data(mem_52_5_W0_data),
    .W0_en(mem_52_5_W0_en),
    .W0_mask(mem_52_5_W0_mask)
  );
  split_mem_0_ext mem_52_6 (
    .R0_addr(mem_52_6_R0_addr),
    .R0_clk(mem_52_6_R0_clk),
    .R0_data(mem_52_6_R0_data),
    .R0_en(mem_52_6_R0_en),
    .W0_addr(mem_52_6_W0_addr),
    .W0_clk(mem_52_6_W0_clk),
    .W0_data(mem_52_6_W0_data),
    .W0_en(mem_52_6_W0_en),
    .W0_mask(mem_52_6_W0_mask)
  );
  split_mem_0_ext mem_52_7 (
    .R0_addr(mem_52_7_R0_addr),
    .R0_clk(mem_52_7_R0_clk),
    .R0_data(mem_52_7_R0_data),
    .R0_en(mem_52_7_R0_en),
    .W0_addr(mem_52_7_W0_addr),
    .W0_clk(mem_52_7_W0_clk),
    .W0_data(mem_52_7_W0_data),
    .W0_en(mem_52_7_W0_en),
    .W0_mask(mem_52_7_W0_mask)
  );
  split_mem_0_ext mem_53_0 (
    .R0_addr(mem_53_0_R0_addr),
    .R0_clk(mem_53_0_R0_clk),
    .R0_data(mem_53_0_R0_data),
    .R0_en(mem_53_0_R0_en),
    .W0_addr(mem_53_0_W0_addr),
    .W0_clk(mem_53_0_W0_clk),
    .W0_data(mem_53_0_W0_data),
    .W0_en(mem_53_0_W0_en),
    .W0_mask(mem_53_0_W0_mask)
  );
  split_mem_0_ext mem_53_1 (
    .R0_addr(mem_53_1_R0_addr),
    .R0_clk(mem_53_1_R0_clk),
    .R0_data(mem_53_1_R0_data),
    .R0_en(mem_53_1_R0_en),
    .W0_addr(mem_53_1_W0_addr),
    .W0_clk(mem_53_1_W0_clk),
    .W0_data(mem_53_1_W0_data),
    .W0_en(mem_53_1_W0_en),
    .W0_mask(mem_53_1_W0_mask)
  );
  split_mem_0_ext mem_53_2 (
    .R0_addr(mem_53_2_R0_addr),
    .R0_clk(mem_53_2_R0_clk),
    .R0_data(mem_53_2_R0_data),
    .R0_en(mem_53_2_R0_en),
    .W0_addr(mem_53_2_W0_addr),
    .W0_clk(mem_53_2_W0_clk),
    .W0_data(mem_53_2_W0_data),
    .W0_en(mem_53_2_W0_en),
    .W0_mask(mem_53_2_W0_mask)
  );
  split_mem_0_ext mem_53_3 (
    .R0_addr(mem_53_3_R0_addr),
    .R0_clk(mem_53_3_R0_clk),
    .R0_data(mem_53_3_R0_data),
    .R0_en(mem_53_3_R0_en),
    .W0_addr(mem_53_3_W0_addr),
    .W0_clk(mem_53_3_W0_clk),
    .W0_data(mem_53_3_W0_data),
    .W0_en(mem_53_3_W0_en),
    .W0_mask(mem_53_3_W0_mask)
  );
  split_mem_0_ext mem_53_4 (
    .R0_addr(mem_53_4_R0_addr),
    .R0_clk(mem_53_4_R0_clk),
    .R0_data(mem_53_4_R0_data),
    .R0_en(mem_53_4_R0_en),
    .W0_addr(mem_53_4_W0_addr),
    .W0_clk(mem_53_4_W0_clk),
    .W0_data(mem_53_4_W0_data),
    .W0_en(mem_53_4_W0_en),
    .W0_mask(mem_53_4_W0_mask)
  );
  split_mem_0_ext mem_53_5 (
    .R0_addr(mem_53_5_R0_addr),
    .R0_clk(mem_53_5_R0_clk),
    .R0_data(mem_53_5_R0_data),
    .R0_en(mem_53_5_R0_en),
    .W0_addr(mem_53_5_W0_addr),
    .W0_clk(mem_53_5_W0_clk),
    .W0_data(mem_53_5_W0_data),
    .W0_en(mem_53_5_W0_en),
    .W0_mask(mem_53_5_W0_mask)
  );
  split_mem_0_ext mem_53_6 (
    .R0_addr(mem_53_6_R0_addr),
    .R0_clk(mem_53_6_R0_clk),
    .R0_data(mem_53_6_R0_data),
    .R0_en(mem_53_6_R0_en),
    .W0_addr(mem_53_6_W0_addr),
    .W0_clk(mem_53_6_W0_clk),
    .W0_data(mem_53_6_W0_data),
    .W0_en(mem_53_6_W0_en),
    .W0_mask(mem_53_6_W0_mask)
  );
  split_mem_0_ext mem_53_7 (
    .R0_addr(mem_53_7_R0_addr),
    .R0_clk(mem_53_7_R0_clk),
    .R0_data(mem_53_7_R0_data),
    .R0_en(mem_53_7_R0_en),
    .W0_addr(mem_53_7_W0_addr),
    .W0_clk(mem_53_7_W0_clk),
    .W0_data(mem_53_7_W0_data),
    .W0_en(mem_53_7_W0_en),
    .W0_mask(mem_53_7_W0_mask)
  );
  split_mem_0_ext mem_54_0 (
    .R0_addr(mem_54_0_R0_addr),
    .R0_clk(mem_54_0_R0_clk),
    .R0_data(mem_54_0_R0_data),
    .R0_en(mem_54_0_R0_en),
    .W0_addr(mem_54_0_W0_addr),
    .W0_clk(mem_54_0_W0_clk),
    .W0_data(mem_54_0_W0_data),
    .W0_en(mem_54_0_W0_en),
    .W0_mask(mem_54_0_W0_mask)
  );
  split_mem_0_ext mem_54_1 (
    .R0_addr(mem_54_1_R0_addr),
    .R0_clk(mem_54_1_R0_clk),
    .R0_data(mem_54_1_R0_data),
    .R0_en(mem_54_1_R0_en),
    .W0_addr(mem_54_1_W0_addr),
    .W0_clk(mem_54_1_W0_clk),
    .W0_data(mem_54_1_W0_data),
    .W0_en(mem_54_1_W0_en),
    .W0_mask(mem_54_1_W0_mask)
  );
  split_mem_0_ext mem_54_2 (
    .R0_addr(mem_54_2_R0_addr),
    .R0_clk(mem_54_2_R0_clk),
    .R0_data(mem_54_2_R0_data),
    .R0_en(mem_54_2_R0_en),
    .W0_addr(mem_54_2_W0_addr),
    .W0_clk(mem_54_2_W0_clk),
    .W0_data(mem_54_2_W0_data),
    .W0_en(mem_54_2_W0_en),
    .W0_mask(mem_54_2_W0_mask)
  );
  split_mem_0_ext mem_54_3 (
    .R0_addr(mem_54_3_R0_addr),
    .R0_clk(mem_54_3_R0_clk),
    .R0_data(mem_54_3_R0_data),
    .R0_en(mem_54_3_R0_en),
    .W0_addr(mem_54_3_W0_addr),
    .W0_clk(mem_54_3_W0_clk),
    .W0_data(mem_54_3_W0_data),
    .W0_en(mem_54_3_W0_en),
    .W0_mask(mem_54_3_W0_mask)
  );
  split_mem_0_ext mem_54_4 (
    .R0_addr(mem_54_4_R0_addr),
    .R0_clk(mem_54_4_R0_clk),
    .R0_data(mem_54_4_R0_data),
    .R0_en(mem_54_4_R0_en),
    .W0_addr(mem_54_4_W0_addr),
    .W0_clk(mem_54_4_W0_clk),
    .W0_data(mem_54_4_W0_data),
    .W0_en(mem_54_4_W0_en),
    .W0_mask(mem_54_4_W0_mask)
  );
  split_mem_0_ext mem_54_5 (
    .R0_addr(mem_54_5_R0_addr),
    .R0_clk(mem_54_5_R0_clk),
    .R0_data(mem_54_5_R0_data),
    .R0_en(mem_54_5_R0_en),
    .W0_addr(mem_54_5_W0_addr),
    .W0_clk(mem_54_5_W0_clk),
    .W0_data(mem_54_5_W0_data),
    .W0_en(mem_54_5_W0_en),
    .W0_mask(mem_54_5_W0_mask)
  );
  split_mem_0_ext mem_54_6 (
    .R0_addr(mem_54_6_R0_addr),
    .R0_clk(mem_54_6_R0_clk),
    .R0_data(mem_54_6_R0_data),
    .R0_en(mem_54_6_R0_en),
    .W0_addr(mem_54_6_W0_addr),
    .W0_clk(mem_54_6_W0_clk),
    .W0_data(mem_54_6_W0_data),
    .W0_en(mem_54_6_W0_en),
    .W0_mask(mem_54_6_W0_mask)
  );
  split_mem_0_ext mem_54_7 (
    .R0_addr(mem_54_7_R0_addr),
    .R0_clk(mem_54_7_R0_clk),
    .R0_data(mem_54_7_R0_data),
    .R0_en(mem_54_7_R0_en),
    .W0_addr(mem_54_7_W0_addr),
    .W0_clk(mem_54_7_W0_clk),
    .W0_data(mem_54_7_W0_data),
    .W0_en(mem_54_7_W0_en),
    .W0_mask(mem_54_7_W0_mask)
  );
  split_mem_0_ext mem_55_0 (
    .R0_addr(mem_55_0_R0_addr),
    .R0_clk(mem_55_0_R0_clk),
    .R0_data(mem_55_0_R0_data),
    .R0_en(mem_55_0_R0_en),
    .W0_addr(mem_55_0_W0_addr),
    .W0_clk(mem_55_0_W0_clk),
    .W0_data(mem_55_0_W0_data),
    .W0_en(mem_55_0_W0_en),
    .W0_mask(mem_55_0_W0_mask)
  );
  split_mem_0_ext mem_55_1 (
    .R0_addr(mem_55_1_R0_addr),
    .R0_clk(mem_55_1_R0_clk),
    .R0_data(mem_55_1_R0_data),
    .R0_en(mem_55_1_R0_en),
    .W0_addr(mem_55_1_W0_addr),
    .W0_clk(mem_55_1_W0_clk),
    .W0_data(mem_55_1_W0_data),
    .W0_en(mem_55_1_W0_en),
    .W0_mask(mem_55_1_W0_mask)
  );
  split_mem_0_ext mem_55_2 (
    .R0_addr(mem_55_2_R0_addr),
    .R0_clk(mem_55_2_R0_clk),
    .R0_data(mem_55_2_R0_data),
    .R0_en(mem_55_2_R0_en),
    .W0_addr(mem_55_2_W0_addr),
    .W0_clk(mem_55_2_W0_clk),
    .W0_data(mem_55_2_W0_data),
    .W0_en(mem_55_2_W0_en),
    .W0_mask(mem_55_2_W0_mask)
  );
  split_mem_0_ext mem_55_3 (
    .R0_addr(mem_55_3_R0_addr),
    .R0_clk(mem_55_3_R0_clk),
    .R0_data(mem_55_3_R0_data),
    .R0_en(mem_55_3_R0_en),
    .W0_addr(mem_55_3_W0_addr),
    .W0_clk(mem_55_3_W0_clk),
    .W0_data(mem_55_3_W0_data),
    .W0_en(mem_55_3_W0_en),
    .W0_mask(mem_55_3_W0_mask)
  );
  split_mem_0_ext mem_55_4 (
    .R0_addr(mem_55_4_R0_addr),
    .R0_clk(mem_55_4_R0_clk),
    .R0_data(mem_55_4_R0_data),
    .R0_en(mem_55_4_R0_en),
    .W0_addr(mem_55_4_W0_addr),
    .W0_clk(mem_55_4_W0_clk),
    .W0_data(mem_55_4_W0_data),
    .W0_en(mem_55_4_W0_en),
    .W0_mask(mem_55_4_W0_mask)
  );
  split_mem_0_ext mem_55_5 (
    .R0_addr(mem_55_5_R0_addr),
    .R0_clk(mem_55_5_R0_clk),
    .R0_data(mem_55_5_R0_data),
    .R0_en(mem_55_5_R0_en),
    .W0_addr(mem_55_5_W0_addr),
    .W0_clk(mem_55_5_W0_clk),
    .W0_data(mem_55_5_W0_data),
    .W0_en(mem_55_5_W0_en),
    .W0_mask(mem_55_5_W0_mask)
  );
  split_mem_0_ext mem_55_6 (
    .R0_addr(mem_55_6_R0_addr),
    .R0_clk(mem_55_6_R0_clk),
    .R0_data(mem_55_6_R0_data),
    .R0_en(mem_55_6_R0_en),
    .W0_addr(mem_55_6_W0_addr),
    .W0_clk(mem_55_6_W0_clk),
    .W0_data(mem_55_6_W0_data),
    .W0_en(mem_55_6_W0_en),
    .W0_mask(mem_55_6_W0_mask)
  );
  split_mem_0_ext mem_55_7 (
    .R0_addr(mem_55_7_R0_addr),
    .R0_clk(mem_55_7_R0_clk),
    .R0_data(mem_55_7_R0_data),
    .R0_en(mem_55_7_R0_en),
    .W0_addr(mem_55_7_W0_addr),
    .W0_clk(mem_55_7_W0_clk),
    .W0_data(mem_55_7_W0_data),
    .W0_en(mem_55_7_W0_en),
    .W0_mask(mem_55_7_W0_mask)
  );
  split_mem_0_ext mem_56_0 (
    .R0_addr(mem_56_0_R0_addr),
    .R0_clk(mem_56_0_R0_clk),
    .R0_data(mem_56_0_R0_data),
    .R0_en(mem_56_0_R0_en),
    .W0_addr(mem_56_0_W0_addr),
    .W0_clk(mem_56_0_W0_clk),
    .W0_data(mem_56_0_W0_data),
    .W0_en(mem_56_0_W0_en),
    .W0_mask(mem_56_0_W0_mask)
  );
  split_mem_0_ext mem_56_1 (
    .R0_addr(mem_56_1_R0_addr),
    .R0_clk(mem_56_1_R0_clk),
    .R0_data(mem_56_1_R0_data),
    .R0_en(mem_56_1_R0_en),
    .W0_addr(mem_56_1_W0_addr),
    .W0_clk(mem_56_1_W0_clk),
    .W0_data(mem_56_1_W0_data),
    .W0_en(mem_56_1_W0_en),
    .W0_mask(mem_56_1_W0_mask)
  );
  split_mem_0_ext mem_56_2 (
    .R0_addr(mem_56_2_R0_addr),
    .R0_clk(mem_56_2_R0_clk),
    .R0_data(mem_56_2_R0_data),
    .R0_en(mem_56_2_R0_en),
    .W0_addr(mem_56_2_W0_addr),
    .W0_clk(mem_56_2_W0_clk),
    .W0_data(mem_56_2_W0_data),
    .W0_en(mem_56_2_W0_en),
    .W0_mask(mem_56_2_W0_mask)
  );
  split_mem_0_ext mem_56_3 (
    .R0_addr(mem_56_3_R0_addr),
    .R0_clk(mem_56_3_R0_clk),
    .R0_data(mem_56_3_R0_data),
    .R0_en(mem_56_3_R0_en),
    .W0_addr(mem_56_3_W0_addr),
    .W0_clk(mem_56_3_W0_clk),
    .W0_data(mem_56_3_W0_data),
    .W0_en(mem_56_3_W0_en),
    .W0_mask(mem_56_3_W0_mask)
  );
  split_mem_0_ext mem_56_4 (
    .R0_addr(mem_56_4_R0_addr),
    .R0_clk(mem_56_4_R0_clk),
    .R0_data(mem_56_4_R0_data),
    .R0_en(mem_56_4_R0_en),
    .W0_addr(mem_56_4_W0_addr),
    .W0_clk(mem_56_4_W0_clk),
    .W0_data(mem_56_4_W0_data),
    .W0_en(mem_56_4_W0_en),
    .W0_mask(mem_56_4_W0_mask)
  );
  split_mem_0_ext mem_56_5 (
    .R0_addr(mem_56_5_R0_addr),
    .R0_clk(mem_56_5_R0_clk),
    .R0_data(mem_56_5_R0_data),
    .R0_en(mem_56_5_R0_en),
    .W0_addr(mem_56_5_W0_addr),
    .W0_clk(mem_56_5_W0_clk),
    .W0_data(mem_56_5_W0_data),
    .W0_en(mem_56_5_W0_en),
    .W0_mask(mem_56_5_W0_mask)
  );
  split_mem_0_ext mem_56_6 (
    .R0_addr(mem_56_6_R0_addr),
    .R0_clk(mem_56_6_R0_clk),
    .R0_data(mem_56_6_R0_data),
    .R0_en(mem_56_6_R0_en),
    .W0_addr(mem_56_6_W0_addr),
    .W0_clk(mem_56_6_W0_clk),
    .W0_data(mem_56_6_W0_data),
    .W0_en(mem_56_6_W0_en),
    .W0_mask(mem_56_6_W0_mask)
  );
  split_mem_0_ext mem_56_7 (
    .R0_addr(mem_56_7_R0_addr),
    .R0_clk(mem_56_7_R0_clk),
    .R0_data(mem_56_7_R0_data),
    .R0_en(mem_56_7_R0_en),
    .W0_addr(mem_56_7_W0_addr),
    .W0_clk(mem_56_7_W0_clk),
    .W0_data(mem_56_7_W0_data),
    .W0_en(mem_56_7_W0_en),
    .W0_mask(mem_56_7_W0_mask)
  );
  split_mem_0_ext mem_57_0 (
    .R0_addr(mem_57_0_R0_addr),
    .R0_clk(mem_57_0_R0_clk),
    .R0_data(mem_57_0_R0_data),
    .R0_en(mem_57_0_R0_en),
    .W0_addr(mem_57_0_W0_addr),
    .W0_clk(mem_57_0_W0_clk),
    .W0_data(mem_57_0_W0_data),
    .W0_en(mem_57_0_W0_en),
    .W0_mask(mem_57_0_W0_mask)
  );
  split_mem_0_ext mem_57_1 (
    .R0_addr(mem_57_1_R0_addr),
    .R0_clk(mem_57_1_R0_clk),
    .R0_data(mem_57_1_R0_data),
    .R0_en(mem_57_1_R0_en),
    .W0_addr(mem_57_1_W0_addr),
    .W0_clk(mem_57_1_W0_clk),
    .W0_data(mem_57_1_W0_data),
    .W0_en(mem_57_1_W0_en),
    .W0_mask(mem_57_1_W0_mask)
  );
  split_mem_0_ext mem_57_2 (
    .R0_addr(mem_57_2_R0_addr),
    .R0_clk(mem_57_2_R0_clk),
    .R0_data(mem_57_2_R0_data),
    .R0_en(mem_57_2_R0_en),
    .W0_addr(mem_57_2_W0_addr),
    .W0_clk(mem_57_2_W0_clk),
    .W0_data(mem_57_2_W0_data),
    .W0_en(mem_57_2_W0_en),
    .W0_mask(mem_57_2_W0_mask)
  );
  split_mem_0_ext mem_57_3 (
    .R0_addr(mem_57_3_R0_addr),
    .R0_clk(mem_57_3_R0_clk),
    .R0_data(mem_57_3_R0_data),
    .R0_en(mem_57_3_R0_en),
    .W0_addr(mem_57_3_W0_addr),
    .W0_clk(mem_57_3_W0_clk),
    .W0_data(mem_57_3_W0_data),
    .W0_en(mem_57_3_W0_en),
    .W0_mask(mem_57_3_W0_mask)
  );
  split_mem_0_ext mem_57_4 (
    .R0_addr(mem_57_4_R0_addr),
    .R0_clk(mem_57_4_R0_clk),
    .R0_data(mem_57_4_R0_data),
    .R0_en(mem_57_4_R0_en),
    .W0_addr(mem_57_4_W0_addr),
    .W0_clk(mem_57_4_W0_clk),
    .W0_data(mem_57_4_W0_data),
    .W0_en(mem_57_4_W0_en),
    .W0_mask(mem_57_4_W0_mask)
  );
  split_mem_0_ext mem_57_5 (
    .R0_addr(mem_57_5_R0_addr),
    .R0_clk(mem_57_5_R0_clk),
    .R0_data(mem_57_5_R0_data),
    .R0_en(mem_57_5_R0_en),
    .W0_addr(mem_57_5_W0_addr),
    .W0_clk(mem_57_5_W0_clk),
    .W0_data(mem_57_5_W0_data),
    .W0_en(mem_57_5_W0_en),
    .W0_mask(mem_57_5_W0_mask)
  );
  split_mem_0_ext mem_57_6 (
    .R0_addr(mem_57_6_R0_addr),
    .R0_clk(mem_57_6_R0_clk),
    .R0_data(mem_57_6_R0_data),
    .R0_en(mem_57_6_R0_en),
    .W0_addr(mem_57_6_W0_addr),
    .W0_clk(mem_57_6_W0_clk),
    .W0_data(mem_57_6_W0_data),
    .W0_en(mem_57_6_W0_en),
    .W0_mask(mem_57_6_W0_mask)
  );
  split_mem_0_ext mem_57_7 (
    .R0_addr(mem_57_7_R0_addr),
    .R0_clk(mem_57_7_R0_clk),
    .R0_data(mem_57_7_R0_data),
    .R0_en(mem_57_7_R0_en),
    .W0_addr(mem_57_7_W0_addr),
    .W0_clk(mem_57_7_W0_clk),
    .W0_data(mem_57_7_W0_data),
    .W0_en(mem_57_7_W0_en),
    .W0_mask(mem_57_7_W0_mask)
  );
  split_mem_0_ext mem_58_0 (
    .R0_addr(mem_58_0_R0_addr),
    .R0_clk(mem_58_0_R0_clk),
    .R0_data(mem_58_0_R0_data),
    .R0_en(mem_58_0_R0_en),
    .W0_addr(mem_58_0_W0_addr),
    .W0_clk(mem_58_0_W0_clk),
    .W0_data(mem_58_0_W0_data),
    .W0_en(mem_58_0_W0_en),
    .W0_mask(mem_58_0_W0_mask)
  );
  split_mem_0_ext mem_58_1 (
    .R0_addr(mem_58_1_R0_addr),
    .R0_clk(mem_58_1_R0_clk),
    .R0_data(mem_58_1_R0_data),
    .R0_en(mem_58_1_R0_en),
    .W0_addr(mem_58_1_W0_addr),
    .W0_clk(mem_58_1_W0_clk),
    .W0_data(mem_58_1_W0_data),
    .W0_en(mem_58_1_W0_en),
    .W0_mask(mem_58_1_W0_mask)
  );
  split_mem_0_ext mem_58_2 (
    .R0_addr(mem_58_2_R0_addr),
    .R0_clk(mem_58_2_R0_clk),
    .R0_data(mem_58_2_R0_data),
    .R0_en(mem_58_2_R0_en),
    .W0_addr(mem_58_2_W0_addr),
    .W0_clk(mem_58_2_W0_clk),
    .W0_data(mem_58_2_W0_data),
    .W0_en(mem_58_2_W0_en),
    .W0_mask(mem_58_2_W0_mask)
  );
  split_mem_0_ext mem_58_3 (
    .R0_addr(mem_58_3_R0_addr),
    .R0_clk(mem_58_3_R0_clk),
    .R0_data(mem_58_3_R0_data),
    .R0_en(mem_58_3_R0_en),
    .W0_addr(mem_58_3_W0_addr),
    .W0_clk(mem_58_3_W0_clk),
    .W0_data(mem_58_3_W0_data),
    .W0_en(mem_58_3_W0_en),
    .W0_mask(mem_58_3_W0_mask)
  );
  split_mem_0_ext mem_58_4 (
    .R0_addr(mem_58_4_R0_addr),
    .R0_clk(mem_58_4_R0_clk),
    .R0_data(mem_58_4_R0_data),
    .R0_en(mem_58_4_R0_en),
    .W0_addr(mem_58_4_W0_addr),
    .W0_clk(mem_58_4_W0_clk),
    .W0_data(mem_58_4_W0_data),
    .W0_en(mem_58_4_W0_en),
    .W0_mask(mem_58_4_W0_mask)
  );
  split_mem_0_ext mem_58_5 (
    .R0_addr(mem_58_5_R0_addr),
    .R0_clk(mem_58_5_R0_clk),
    .R0_data(mem_58_5_R0_data),
    .R0_en(mem_58_5_R0_en),
    .W0_addr(mem_58_5_W0_addr),
    .W0_clk(mem_58_5_W0_clk),
    .W0_data(mem_58_5_W0_data),
    .W0_en(mem_58_5_W0_en),
    .W0_mask(mem_58_5_W0_mask)
  );
  split_mem_0_ext mem_58_6 (
    .R0_addr(mem_58_6_R0_addr),
    .R0_clk(mem_58_6_R0_clk),
    .R0_data(mem_58_6_R0_data),
    .R0_en(mem_58_6_R0_en),
    .W0_addr(mem_58_6_W0_addr),
    .W0_clk(mem_58_6_W0_clk),
    .W0_data(mem_58_6_W0_data),
    .W0_en(mem_58_6_W0_en),
    .W0_mask(mem_58_6_W0_mask)
  );
  split_mem_0_ext mem_58_7 (
    .R0_addr(mem_58_7_R0_addr),
    .R0_clk(mem_58_7_R0_clk),
    .R0_data(mem_58_7_R0_data),
    .R0_en(mem_58_7_R0_en),
    .W0_addr(mem_58_7_W0_addr),
    .W0_clk(mem_58_7_W0_clk),
    .W0_data(mem_58_7_W0_data),
    .W0_en(mem_58_7_W0_en),
    .W0_mask(mem_58_7_W0_mask)
  );
  split_mem_0_ext mem_59_0 (
    .R0_addr(mem_59_0_R0_addr),
    .R0_clk(mem_59_0_R0_clk),
    .R0_data(mem_59_0_R0_data),
    .R0_en(mem_59_0_R0_en),
    .W0_addr(mem_59_0_W0_addr),
    .W0_clk(mem_59_0_W0_clk),
    .W0_data(mem_59_0_W0_data),
    .W0_en(mem_59_0_W0_en),
    .W0_mask(mem_59_0_W0_mask)
  );
  split_mem_0_ext mem_59_1 (
    .R0_addr(mem_59_1_R0_addr),
    .R0_clk(mem_59_1_R0_clk),
    .R0_data(mem_59_1_R0_data),
    .R0_en(mem_59_1_R0_en),
    .W0_addr(mem_59_1_W0_addr),
    .W0_clk(mem_59_1_W0_clk),
    .W0_data(mem_59_1_W0_data),
    .W0_en(mem_59_1_W0_en),
    .W0_mask(mem_59_1_W0_mask)
  );
  split_mem_0_ext mem_59_2 (
    .R0_addr(mem_59_2_R0_addr),
    .R0_clk(mem_59_2_R0_clk),
    .R0_data(mem_59_2_R0_data),
    .R0_en(mem_59_2_R0_en),
    .W0_addr(mem_59_2_W0_addr),
    .W0_clk(mem_59_2_W0_clk),
    .W0_data(mem_59_2_W0_data),
    .W0_en(mem_59_2_W0_en),
    .W0_mask(mem_59_2_W0_mask)
  );
  split_mem_0_ext mem_59_3 (
    .R0_addr(mem_59_3_R0_addr),
    .R0_clk(mem_59_3_R0_clk),
    .R0_data(mem_59_3_R0_data),
    .R0_en(mem_59_3_R0_en),
    .W0_addr(mem_59_3_W0_addr),
    .W0_clk(mem_59_3_W0_clk),
    .W0_data(mem_59_3_W0_data),
    .W0_en(mem_59_3_W0_en),
    .W0_mask(mem_59_3_W0_mask)
  );
  split_mem_0_ext mem_59_4 (
    .R0_addr(mem_59_4_R0_addr),
    .R0_clk(mem_59_4_R0_clk),
    .R0_data(mem_59_4_R0_data),
    .R0_en(mem_59_4_R0_en),
    .W0_addr(mem_59_4_W0_addr),
    .W0_clk(mem_59_4_W0_clk),
    .W0_data(mem_59_4_W0_data),
    .W0_en(mem_59_4_W0_en),
    .W0_mask(mem_59_4_W0_mask)
  );
  split_mem_0_ext mem_59_5 (
    .R0_addr(mem_59_5_R0_addr),
    .R0_clk(mem_59_5_R0_clk),
    .R0_data(mem_59_5_R0_data),
    .R0_en(mem_59_5_R0_en),
    .W0_addr(mem_59_5_W0_addr),
    .W0_clk(mem_59_5_W0_clk),
    .W0_data(mem_59_5_W0_data),
    .W0_en(mem_59_5_W0_en),
    .W0_mask(mem_59_5_W0_mask)
  );
  split_mem_0_ext mem_59_6 (
    .R0_addr(mem_59_6_R0_addr),
    .R0_clk(mem_59_6_R0_clk),
    .R0_data(mem_59_6_R0_data),
    .R0_en(mem_59_6_R0_en),
    .W0_addr(mem_59_6_W0_addr),
    .W0_clk(mem_59_6_W0_clk),
    .W0_data(mem_59_6_W0_data),
    .W0_en(mem_59_6_W0_en),
    .W0_mask(mem_59_6_W0_mask)
  );
  split_mem_0_ext mem_59_7 (
    .R0_addr(mem_59_7_R0_addr),
    .R0_clk(mem_59_7_R0_clk),
    .R0_data(mem_59_7_R0_data),
    .R0_en(mem_59_7_R0_en),
    .W0_addr(mem_59_7_W0_addr),
    .W0_clk(mem_59_7_W0_clk),
    .W0_data(mem_59_7_W0_data),
    .W0_en(mem_59_7_W0_en),
    .W0_mask(mem_59_7_W0_mask)
  );
  split_mem_0_ext mem_60_0 (
    .R0_addr(mem_60_0_R0_addr),
    .R0_clk(mem_60_0_R0_clk),
    .R0_data(mem_60_0_R0_data),
    .R0_en(mem_60_0_R0_en),
    .W0_addr(mem_60_0_W0_addr),
    .W0_clk(mem_60_0_W0_clk),
    .W0_data(mem_60_0_W0_data),
    .W0_en(mem_60_0_W0_en),
    .W0_mask(mem_60_0_W0_mask)
  );
  split_mem_0_ext mem_60_1 (
    .R0_addr(mem_60_1_R0_addr),
    .R0_clk(mem_60_1_R0_clk),
    .R0_data(mem_60_1_R0_data),
    .R0_en(mem_60_1_R0_en),
    .W0_addr(mem_60_1_W0_addr),
    .W0_clk(mem_60_1_W0_clk),
    .W0_data(mem_60_1_W0_data),
    .W0_en(mem_60_1_W0_en),
    .W0_mask(mem_60_1_W0_mask)
  );
  split_mem_0_ext mem_60_2 (
    .R0_addr(mem_60_2_R0_addr),
    .R0_clk(mem_60_2_R0_clk),
    .R0_data(mem_60_2_R0_data),
    .R0_en(mem_60_2_R0_en),
    .W0_addr(mem_60_2_W0_addr),
    .W0_clk(mem_60_2_W0_clk),
    .W0_data(mem_60_2_W0_data),
    .W0_en(mem_60_2_W0_en),
    .W0_mask(mem_60_2_W0_mask)
  );
  split_mem_0_ext mem_60_3 (
    .R0_addr(mem_60_3_R0_addr),
    .R0_clk(mem_60_3_R0_clk),
    .R0_data(mem_60_3_R0_data),
    .R0_en(mem_60_3_R0_en),
    .W0_addr(mem_60_3_W0_addr),
    .W0_clk(mem_60_3_W0_clk),
    .W0_data(mem_60_3_W0_data),
    .W0_en(mem_60_3_W0_en),
    .W0_mask(mem_60_3_W0_mask)
  );
  split_mem_0_ext mem_60_4 (
    .R0_addr(mem_60_4_R0_addr),
    .R0_clk(mem_60_4_R0_clk),
    .R0_data(mem_60_4_R0_data),
    .R0_en(mem_60_4_R0_en),
    .W0_addr(mem_60_4_W0_addr),
    .W0_clk(mem_60_4_W0_clk),
    .W0_data(mem_60_4_W0_data),
    .W0_en(mem_60_4_W0_en),
    .W0_mask(mem_60_4_W0_mask)
  );
  split_mem_0_ext mem_60_5 (
    .R0_addr(mem_60_5_R0_addr),
    .R0_clk(mem_60_5_R0_clk),
    .R0_data(mem_60_5_R0_data),
    .R0_en(mem_60_5_R0_en),
    .W0_addr(mem_60_5_W0_addr),
    .W0_clk(mem_60_5_W0_clk),
    .W0_data(mem_60_5_W0_data),
    .W0_en(mem_60_5_W0_en),
    .W0_mask(mem_60_5_W0_mask)
  );
  split_mem_0_ext mem_60_6 (
    .R0_addr(mem_60_6_R0_addr),
    .R0_clk(mem_60_6_R0_clk),
    .R0_data(mem_60_6_R0_data),
    .R0_en(mem_60_6_R0_en),
    .W0_addr(mem_60_6_W0_addr),
    .W0_clk(mem_60_6_W0_clk),
    .W0_data(mem_60_6_W0_data),
    .W0_en(mem_60_6_W0_en),
    .W0_mask(mem_60_6_W0_mask)
  );
  split_mem_0_ext mem_60_7 (
    .R0_addr(mem_60_7_R0_addr),
    .R0_clk(mem_60_7_R0_clk),
    .R0_data(mem_60_7_R0_data),
    .R0_en(mem_60_7_R0_en),
    .W0_addr(mem_60_7_W0_addr),
    .W0_clk(mem_60_7_W0_clk),
    .W0_data(mem_60_7_W0_data),
    .W0_en(mem_60_7_W0_en),
    .W0_mask(mem_60_7_W0_mask)
  );
  split_mem_0_ext mem_61_0 (
    .R0_addr(mem_61_0_R0_addr),
    .R0_clk(mem_61_0_R0_clk),
    .R0_data(mem_61_0_R0_data),
    .R0_en(mem_61_0_R0_en),
    .W0_addr(mem_61_0_W0_addr),
    .W0_clk(mem_61_0_W0_clk),
    .W0_data(mem_61_0_W0_data),
    .W0_en(mem_61_0_W0_en),
    .W0_mask(mem_61_0_W0_mask)
  );
  split_mem_0_ext mem_61_1 (
    .R0_addr(mem_61_1_R0_addr),
    .R0_clk(mem_61_1_R0_clk),
    .R0_data(mem_61_1_R0_data),
    .R0_en(mem_61_1_R0_en),
    .W0_addr(mem_61_1_W0_addr),
    .W0_clk(mem_61_1_W0_clk),
    .W0_data(mem_61_1_W0_data),
    .W0_en(mem_61_1_W0_en),
    .W0_mask(mem_61_1_W0_mask)
  );
  split_mem_0_ext mem_61_2 (
    .R0_addr(mem_61_2_R0_addr),
    .R0_clk(mem_61_2_R0_clk),
    .R0_data(mem_61_2_R0_data),
    .R0_en(mem_61_2_R0_en),
    .W0_addr(mem_61_2_W0_addr),
    .W0_clk(mem_61_2_W0_clk),
    .W0_data(mem_61_2_W0_data),
    .W0_en(mem_61_2_W0_en),
    .W0_mask(mem_61_2_W0_mask)
  );
  split_mem_0_ext mem_61_3 (
    .R0_addr(mem_61_3_R0_addr),
    .R0_clk(mem_61_3_R0_clk),
    .R0_data(mem_61_3_R0_data),
    .R0_en(mem_61_3_R0_en),
    .W0_addr(mem_61_3_W0_addr),
    .W0_clk(mem_61_3_W0_clk),
    .W0_data(mem_61_3_W0_data),
    .W0_en(mem_61_3_W0_en),
    .W0_mask(mem_61_3_W0_mask)
  );
  split_mem_0_ext mem_61_4 (
    .R0_addr(mem_61_4_R0_addr),
    .R0_clk(mem_61_4_R0_clk),
    .R0_data(mem_61_4_R0_data),
    .R0_en(mem_61_4_R0_en),
    .W0_addr(mem_61_4_W0_addr),
    .W0_clk(mem_61_4_W0_clk),
    .W0_data(mem_61_4_W0_data),
    .W0_en(mem_61_4_W0_en),
    .W0_mask(mem_61_4_W0_mask)
  );
  split_mem_0_ext mem_61_5 (
    .R0_addr(mem_61_5_R0_addr),
    .R0_clk(mem_61_5_R0_clk),
    .R0_data(mem_61_5_R0_data),
    .R0_en(mem_61_5_R0_en),
    .W0_addr(mem_61_5_W0_addr),
    .W0_clk(mem_61_5_W0_clk),
    .W0_data(mem_61_5_W0_data),
    .W0_en(mem_61_5_W0_en),
    .W0_mask(mem_61_5_W0_mask)
  );
  split_mem_0_ext mem_61_6 (
    .R0_addr(mem_61_6_R0_addr),
    .R0_clk(mem_61_6_R0_clk),
    .R0_data(mem_61_6_R0_data),
    .R0_en(mem_61_6_R0_en),
    .W0_addr(mem_61_6_W0_addr),
    .W0_clk(mem_61_6_W0_clk),
    .W0_data(mem_61_6_W0_data),
    .W0_en(mem_61_6_W0_en),
    .W0_mask(mem_61_6_W0_mask)
  );
  split_mem_0_ext mem_61_7 (
    .R0_addr(mem_61_7_R0_addr),
    .R0_clk(mem_61_7_R0_clk),
    .R0_data(mem_61_7_R0_data),
    .R0_en(mem_61_7_R0_en),
    .W0_addr(mem_61_7_W0_addr),
    .W0_clk(mem_61_7_W0_clk),
    .W0_data(mem_61_7_W0_data),
    .W0_en(mem_61_7_W0_en),
    .W0_mask(mem_61_7_W0_mask)
  );
  split_mem_0_ext mem_62_0 (
    .R0_addr(mem_62_0_R0_addr),
    .R0_clk(mem_62_0_R0_clk),
    .R0_data(mem_62_0_R0_data),
    .R0_en(mem_62_0_R0_en),
    .W0_addr(mem_62_0_W0_addr),
    .W0_clk(mem_62_0_W0_clk),
    .W0_data(mem_62_0_W0_data),
    .W0_en(mem_62_0_W0_en),
    .W0_mask(mem_62_0_W0_mask)
  );
  split_mem_0_ext mem_62_1 (
    .R0_addr(mem_62_1_R0_addr),
    .R0_clk(mem_62_1_R0_clk),
    .R0_data(mem_62_1_R0_data),
    .R0_en(mem_62_1_R0_en),
    .W0_addr(mem_62_1_W0_addr),
    .W0_clk(mem_62_1_W0_clk),
    .W0_data(mem_62_1_W0_data),
    .W0_en(mem_62_1_W0_en),
    .W0_mask(mem_62_1_W0_mask)
  );
  split_mem_0_ext mem_62_2 (
    .R0_addr(mem_62_2_R0_addr),
    .R0_clk(mem_62_2_R0_clk),
    .R0_data(mem_62_2_R0_data),
    .R0_en(mem_62_2_R0_en),
    .W0_addr(mem_62_2_W0_addr),
    .W0_clk(mem_62_2_W0_clk),
    .W0_data(mem_62_2_W0_data),
    .W0_en(mem_62_2_W0_en),
    .W0_mask(mem_62_2_W0_mask)
  );
  split_mem_0_ext mem_62_3 (
    .R0_addr(mem_62_3_R0_addr),
    .R0_clk(mem_62_3_R0_clk),
    .R0_data(mem_62_3_R0_data),
    .R0_en(mem_62_3_R0_en),
    .W0_addr(mem_62_3_W0_addr),
    .W0_clk(mem_62_3_W0_clk),
    .W0_data(mem_62_3_W0_data),
    .W0_en(mem_62_3_W0_en),
    .W0_mask(mem_62_3_W0_mask)
  );
  split_mem_0_ext mem_62_4 (
    .R0_addr(mem_62_4_R0_addr),
    .R0_clk(mem_62_4_R0_clk),
    .R0_data(mem_62_4_R0_data),
    .R0_en(mem_62_4_R0_en),
    .W0_addr(mem_62_4_W0_addr),
    .W0_clk(mem_62_4_W0_clk),
    .W0_data(mem_62_4_W0_data),
    .W0_en(mem_62_4_W0_en),
    .W0_mask(mem_62_4_W0_mask)
  );
  split_mem_0_ext mem_62_5 (
    .R0_addr(mem_62_5_R0_addr),
    .R0_clk(mem_62_5_R0_clk),
    .R0_data(mem_62_5_R0_data),
    .R0_en(mem_62_5_R0_en),
    .W0_addr(mem_62_5_W0_addr),
    .W0_clk(mem_62_5_W0_clk),
    .W0_data(mem_62_5_W0_data),
    .W0_en(mem_62_5_W0_en),
    .W0_mask(mem_62_5_W0_mask)
  );
  split_mem_0_ext mem_62_6 (
    .R0_addr(mem_62_6_R0_addr),
    .R0_clk(mem_62_6_R0_clk),
    .R0_data(mem_62_6_R0_data),
    .R0_en(mem_62_6_R0_en),
    .W0_addr(mem_62_6_W0_addr),
    .W0_clk(mem_62_6_W0_clk),
    .W0_data(mem_62_6_W0_data),
    .W0_en(mem_62_6_W0_en),
    .W0_mask(mem_62_6_W0_mask)
  );
  split_mem_0_ext mem_62_7 (
    .R0_addr(mem_62_7_R0_addr),
    .R0_clk(mem_62_7_R0_clk),
    .R0_data(mem_62_7_R0_data),
    .R0_en(mem_62_7_R0_en),
    .W0_addr(mem_62_7_W0_addr),
    .W0_clk(mem_62_7_W0_clk),
    .W0_data(mem_62_7_W0_data),
    .W0_en(mem_62_7_W0_en),
    .W0_mask(mem_62_7_W0_mask)
  );
  split_mem_0_ext mem_63_0 (
    .R0_addr(mem_63_0_R0_addr),
    .R0_clk(mem_63_0_R0_clk),
    .R0_data(mem_63_0_R0_data),
    .R0_en(mem_63_0_R0_en),
    .W0_addr(mem_63_0_W0_addr),
    .W0_clk(mem_63_0_W0_clk),
    .W0_data(mem_63_0_W0_data),
    .W0_en(mem_63_0_W0_en),
    .W0_mask(mem_63_0_W0_mask)
  );
  split_mem_0_ext mem_63_1 (
    .R0_addr(mem_63_1_R0_addr),
    .R0_clk(mem_63_1_R0_clk),
    .R0_data(mem_63_1_R0_data),
    .R0_en(mem_63_1_R0_en),
    .W0_addr(mem_63_1_W0_addr),
    .W0_clk(mem_63_1_W0_clk),
    .W0_data(mem_63_1_W0_data),
    .W0_en(mem_63_1_W0_en),
    .W0_mask(mem_63_1_W0_mask)
  );
  split_mem_0_ext mem_63_2 (
    .R0_addr(mem_63_2_R0_addr),
    .R0_clk(mem_63_2_R0_clk),
    .R0_data(mem_63_2_R0_data),
    .R0_en(mem_63_2_R0_en),
    .W0_addr(mem_63_2_W0_addr),
    .W0_clk(mem_63_2_W0_clk),
    .W0_data(mem_63_2_W0_data),
    .W0_en(mem_63_2_W0_en),
    .W0_mask(mem_63_2_W0_mask)
  );
  split_mem_0_ext mem_63_3 (
    .R0_addr(mem_63_3_R0_addr),
    .R0_clk(mem_63_3_R0_clk),
    .R0_data(mem_63_3_R0_data),
    .R0_en(mem_63_3_R0_en),
    .W0_addr(mem_63_3_W0_addr),
    .W0_clk(mem_63_3_W0_clk),
    .W0_data(mem_63_3_W0_data),
    .W0_en(mem_63_3_W0_en),
    .W0_mask(mem_63_3_W0_mask)
  );
  split_mem_0_ext mem_63_4 (
    .R0_addr(mem_63_4_R0_addr),
    .R0_clk(mem_63_4_R0_clk),
    .R0_data(mem_63_4_R0_data),
    .R0_en(mem_63_4_R0_en),
    .W0_addr(mem_63_4_W0_addr),
    .W0_clk(mem_63_4_W0_clk),
    .W0_data(mem_63_4_W0_data),
    .W0_en(mem_63_4_W0_en),
    .W0_mask(mem_63_4_W0_mask)
  );
  split_mem_0_ext mem_63_5 (
    .R0_addr(mem_63_5_R0_addr),
    .R0_clk(mem_63_5_R0_clk),
    .R0_data(mem_63_5_R0_data),
    .R0_en(mem_63_5_R0_en),
    .W0_addr(mem_63_5_W0_addr),
    .W0_clk(mem_63_5_W0_clk),
    .W0_data(mem_63_5_W0_data),
    .W0_en(mem_63_5_W0_en),
    .W0_mask(mem_63_5_W0_mask)
  );
  split_mem_0_ext mem_63_6 (
    .R0_addr(mem_63_6_R0_addr),
    .R0_clk(mem_63_6_R0_clk),
    .R0_data(mem_63_6_R0_data),
    .R0_en(mem_63_6_R0_en),
    .W0_addr(mem_63_6_W0_addr),
    .W0_clk(mem_63_6_W0_clk),
    .W0_data(mem_63_6_W0_data),
    .W0_en(mem_63_6_W0_en),
    .W0_mask(mem_63_6_W0_mask)
  );
  split_mem_0_ext mem_63_7 (
    .R0_addr(mem_63_7_R0_addr),
    .R0_clk(mem_63_7_R0_clk),
    .R0_data(mem_63_7_R0_data),
    .R0_en(mem_63_7_R0_en),
    .W0_addr(mem_63_7_W0_addr),
    .W0_clk(mem_63_7_W0_clk),
    .W0_data(mem_63_7_W0_data),
    .W0_en(mem_63_7_W0_en),
    .W0_mask(mem_63_7_W0_mask)
  );
  split_mem_0_ext mem_64_0 (
    .R0_addr(mem_64_0_R0_addr),
    .R0_clk(mem_64_0_R0_clk),
    .R0_data(mem_64_0_R0_data),
    .R0_en(mem_64_0_R0_en),
    .W0_addr(mem_64_0_W0_addr),
    .W0_clk(mem_64_0_W0_clk),
    .W0_data(mem_64_0_W0_data),
    .W0_en(mem_64_0_W0_en),
    .W0_mask(mem_64_0_W0_mask)
  );
  split_mem_0_ext mem_64_1 (
    .R0_addr(mem_64_1_R0_addr),
    .R0_clk(mem_64_1_R0_clk),
    .R0_data(mem_64_1_R0_data),
    .R0_en(mem_64_1_R0_en),
    .W0_addr(mem_64_1_W0_addr),
    .W0_clk(mem_64_1_W0_clk),
    .W0_data(mem_64_1_W0_data),
    .W0_en(mem_64_1_W0_en),
    .W0_mask(mem_64_1_W0_mask)
  );
  split_mem_0_ext mem_64_2 (
    .R0_addr(mem_64_2_R0_addr),
    .R0_clk(mem_64_2_R0_clk),
    .R0_data(mem_64_2_R0_data),
    .R0_en(mem_64_2_R0_en),
    .W0_addr(mem_64_2_W0_addr),
    .W0_clk(mem_64_2_W0_clk),
    .W0_data(mem_64_2_W0_data),
    .W0_en(mem_64_2_W0_en),
    .W0_mask(mem_64_2_W0_mask)
  );
  split_mem_0_ext mem_64_3 (
    .R0_addr(mem_64_3_R0_addr),
    .R0_clk(mem_64_3_R0_clk),
    .R0_data(mem_64_3_R0_data),
    .R0_en(mem_64_3_R0_en),
    .W0_addr(mem_64_3_W0_addr),
    .W0_clk(mem_64_3_W0_clk),
    .W0_data(mem_64_3_W0_data),
    .W0_en(mem_64_3_W0_en),
    .W0_mask(mem_64_3_W0_mask)
  );
  split_mem_0_ext mem_64_4 (
    .R0_addr(mem_64_4_R0_addr),
    .R0_clk(mem_64_4_R0_clk),
    .R0_data(mem_64_4_R0_data),
    .R0_en(mem_64_4_R0_en),
    .W0_addr(mem_64_4_W0_addr),
    .W0_clk(mem_64_4_W0_clk),
    .W0_data(mem_64_4_W0_data),
    .W0_en(mem_64_4_W0_en),
    .W0_mask(mem_64_4_W0_mask)
  );
  split_mem_0_ext mem_64_5 (
    .R0_addr(mem_64_5_R0_addr),
    .R0_clk(mem_64_5_R0_clk),
    .R0_data(mem_64_5_R0_data),
    .R0_en(mem_64_5_R0_en),
    .W0_addr(mem_64_5_W0_addr),
    .W0_clk(mem_64_5_W0_clk),
    .W0_data(mem_64_5_W0_data),
    .W0_en(mem_64_5_W0_en),
    .W0_mask(mem_64_5_W0_mask)
  );
  split_mem_0_ext mem_64_6 (
    .R0_addr(mem_64_6_R0_addr),
    .R0_clk(mem_64_6_R0_clk),
    .R0_data(mem_64_6_R0_data),
    .R0_en(mem_64_6_R0_en),
    .W0_addr(mem_64_6_W0_addr),
    .W0_clk(mem_64_6_W0_clk),
    .W0_data(mem_64_6_W0_data),
    .W0_en(mem_64_6_W0_en),
    .W0_mask(mem_64_6_W0_mask)
  );
  split_mem_0_ext mem_64_7 (
    .R0_addr(mem_64_7_R0_addr),
    .R0_clk(mem_64_7_R0_clk),
    .R0_data(mem_64_7_R0_data),
    .R0_en(mem_64_7_R0_en),
    .W0_addr(mem_64_7_W0_addr),
    .W0_clk(mem_64_7_W0_clk),
    .W0_data(mem_64_7_W0_data),
    .W0_en(mem_64_7_W0_en),
    .W0_mask(mem_64_7_W0_mask)
  );
  split_mem_0_ext mem_65_0 (
    .R0_addr(mem_65_0_R0_addr),
    .R0_clk(mem_65_0_R0_clk),
    .R0_data(mem_65_0_R0_data),
    .R0_en(mem_65_0_R0_en),
    .W0_addr(mem_65_0_W0_addr),
    .W0_clk(mem_65_0_W0_clk),
    .W0_data(mem_65_0_W0_data),
    .W0_en(mem_65_0_W0_en),
    .W0_mask(mem_65_0_W0_mask)
  );
  split_mem_0_ext mem_65_1 (
    .R0_addr(mem_65_1_R0_addr),
    .R0_clk(mem_65_1_R0_clk),
    .R0_data(mem_65_1_R0_data),
    .R0_en(mem_65_1_R0_en),
    .W0_addr(mem_65_1_W0_addr),
    .W0_clk(mem_65_1_W0_clk),
    .W0_data(mem_65_1_W0_data),
    .W0_en(mem_65_1_W0_en),
    .W0_mask(mem_65_1_W0_mask)
  );
  split_mem_0_ext mem_65_2 (
    .R0_addr(mem_65_2_R0_addr),
    .R0_clk(mem_65_2_R0_clk),
    .R0_data(mem_65_2_R0_data),
    .R0_en(mem_65_2_R0_en),
    .W0_addr(mem_65_2_W0_addr),
    .W0_clk(mem_65_2_W0_clk),
    .W0_data(mem_65_2_W0_data),
    .W0_en(mem_65_2_W0_en),
    .W0_mask(mem_65_2_W0_mask)
  );
  split_mem_0_ext mem_65_3 (
    .R0_addr(mem_65_3_R0_addr),
    .R0_clk(mem_65_3_R0_clk),
    .R0_data(mem_65_3_R0_data),
    .R0_en(mem_65_3_R0_en),
    .W0_addr(mem_65_3_W0_addr),
    .W0_clk(mem_65_3_W0_clk),
    .W0_data(mem_65_3_W0_data),
    .W0_en(mem_65_3_W0_en),
    .W0_mask(mem_65_3_W0_mask)
  );
  split_mem_0_ext mem_65_4 (
    .R0_addr(mem_65_4_R0_addr),
    .R0_clk(mem_65_4_R0_clk),
    .R0_data(mem_65_4_R0_data),
    .R0_en(mem_65_4_R0_en),
    .W0_addr(mem_65_4_W0_addr),
    .W0_clk(mem_65_4_W0_clk),
    .W0_data(mem_65_4_W0_data),
    .W0_en(mem_65_4_W0_en),
    .W0_mask(mem_65_4_W0_mask)
  );
  split_mem_0_ext mem_65_5 (
    .R0_addr(mem_65_5_R0_addr),
    .R0_clk(mem_65_5_R0_clk),
    .R0_data(mem_65_5_R0_data),
    .R0_en(mem_65_5_R0_en),
    .W0_addr(mem_65_5_W0_addr),
    .W0_clk(mem_65_5_W0_clk),
    .W0_data(mem_65_5_W0_data),
    .W0_en(mem_65_5_W0_en),
    .W0_mask(mem_65_5_W0_mask)
  );
  split_mem_0_ext mem_65_6 (
    .R0_addr(mem_65_6_R0_addr),
    .R0_clk(mem_65_6_R0_clk),
    .R0_data(mem_65_6_R0_data),
    .R0_en(mem_65_6_R0_en),
    .W0_addr(mem_65_6_W0_addr),
    .W0_clk(mem_65_6_W0_clk),
    .W0_data(mem_65_6_W0_data),
    .W0_en(mem_65_6_W0_en),
    .W0_mask(mem_65_6_W0_mask)
  );
  split_mem_0_ext mem_65_7 (
    .R0_addr(mem_65_7_R0_addr),
    .R0_clk(mem_65_7_R0_clk),
    .R0_data(mem_65_7_R0_data),
    .R0_en(mem_65_7_R0_en),
    .W0_addr(mem_65_7_W0_addr),
    .W0_clk(mem_65_7_W0_clk),
    .W0_data(mem_65_7_W0_data),
    .W0_en(mem_65_7_W0_en),
    .W0_mask(mem_65_7_W0_mask)
  );
  split_mem_0_ext mem_66_0 (
    .R0_addr(mem_66_0_R0_addr),
    .R0_clk(mem_66_0_R0_clk),
    .R0_data(mem_66_0_R0_data),
    .R0_en(mem_66_0_R0_en),
    .W0_addr(mem_66_0_W0_addr),
    .W0_clk(mem_66_0_W0_clk),
    .W0_data(mem_66_0_W0_data),
    .W0_en(mem_66_0_W0_en),
    .W0_mask(mem_66_0_W0_mask)
  );
  split_mem_0_ext mem_66_1 (
    .R0_addr(mem_66_1_R0_addr),
    .R0_clk(mem_66_1_R0_clk),
    .R0_data(mem_66_1_R0_data),
    .R0_en(mem_66_1_R0_en),
    .W0_addr(mem_66_1_W0_addr),
    .W0_clk(mem_66_1_W0_clk),
    .W0_data(mem_66_1_W0_data),
    .W0_en(mem_66_1_W0_en),
    .W0_mask(mem_66_1_W0_mask)
  );
  split_mem_0_ext mem_66_2 (
    .R0_addr(mem_66_2_R0_addr),
    .R0_clk(mem_66_2_R0_clk),
    .R0_data(mem_66_2_R0_data),
    .R0_en(mem_66_2_R0_en),
    .W0_addr(mem_66_2_W0_addr),
    .W0_clk(mem_66_2_W0_clk),
    .W0_data(mem_66_2_W0_data),
    .W0_en(mem_66_2_W0_en),
    .W0_mask(mem_66_2_W0_mask)
  );
  split_mem_0_ext mem_66_3 (
    .R0_addr(mem_66_3_R0_addr),
    .R0_clk(mem_66_3_R0_clk),
    .R0_data(mem_66_3_R0_data),
    .R0_en(mem_66_3_R0_en),
    .W0_addr(mem_66_3_W0_addr),
    .W0_clk(mem_66_3_W0_clk),
    .W0_data(mem_66_3_W0_data),
    .W0_en(mem_66_3_W0_en),
    .W0_mask(mem_66_3_W0_mask)
  );
  split_mem_0_ext mem_66_4 (
    .R0_addr(mem_66_4_R0_addr),
    .R0_clk(mem_66_4_R0_clk),
    .R0_data(mem_66_4_R0_data),
    .R0_en(mem_66_4_R0_en),
    .W0_addr(mem_66_4_W0_addr),
    .W0_clk(mem_66_4_W0_clk),
    .W0_data(mem_66_4_W0_data),
    .W0_en(mem_66_4_W0_en),
    .W0_mask(mem_66_4_W0_mask)
  );
  split_mem_0_ext mem_66_5 (
    .R0_addr(mem_66_5_R0_addr),
    .R0_clk(mem_66_5_R0_clk),
    .R0_data(mem_66_5_R0_data),
    .R0_en(mem_66_5_R0_en),
    .W0_addr(mem_66_5_W0_addr),
    .W0_clk(mem_66_5_W0_clk),
    .W0_data(mem_66_5_W0_data),
    .W0_en(mem_66_5_W0_en),
    .W0_mask(mem_66_5_W0_mask)
  );
  split_mem_0_ext mem_66_6 (
    .R0_addr(mem_66_6_R0_addr),
    .R0_clk(mem_66_6_R0_clk),
    .R0_data(mem_66_6_R0_data),
    .R0_en(mem_66_6_R0_en),
    .W0_addr(mem_66_6_W0_addr),
    .W0_clk(mem_66_6_W0_clk),
    .W0_data(mem_66_6_W0_data),
    .W0_en(mem_66_6_W0_en),
    .W0_mask(mem_66_6_W0_mask)
  );
  split_mem_0_ext mem_66_7 (
    .R0_addr(mem_66_7_R0_addr),
    .R0_clk(mem_66_7_R0_clk),
    .R0_data(mem_66_7_R0_data),
    .R0_en(mem_66_7_R0_en),
    .W0_addr(mem_66_7_W0_addr),
    .W0_clk(mem_66_7_W0_clk),
    .W0_data(mem_66_7_W0_data),
    .W0_en(mem_66_7_W0_en),
    .W0_mask(mem_66_7_W0_mask)
  );
  split_mem_0_ext mem_67_0 (
    .R0_addr(mem_67_0_R0_addr),
    .R0_clk(mem_67_0_R0_clk),
    .R0_data(mem_67_0_R0_data),
    .R0_en(mem_67_0_R0_en),
    .W0_addr(mem_67_0_W0_addr),
    .W0_clk(mem_67_0_W0_clk),
    .W0_data(mem_67_0_W0_data),
    .W0_en(mem_67_0_W0_en),
    .W0_mask(mem_67_0_W0_mask)
  );
  split_mem_0_ext mem_67_1 (
    .R0_addr(mem_67_1_R0_addr),
    .R0_clk(mem_67_1_R0_clk),
    .R0_data(mem_67_1_R0_data),
    .R0_en(mem_67_1_R0_en),
    .W0_addr(mem_67_1_W0_addr),
    .W0_clk(mem_67_1_W0_clk),
    .W0_data(mem_67_1_W0_data),
    .W0_en(mem_67_1_W0_en),
    .W0_mask(mem_67_1_W0_mask)
  );
  split_mem_0_ext mem_67_2 (
    .R0_addr(mem_67_2_R0_addr),
    .R0_clk(mem_67_2_R0_clk),
    .R0_data(mem_67_2_R0_data),
    .R0_en(mem_67_2_R0_en),
    .W0_addr(mem_67_2_W0_addr),
    .W0_clk(mem_67_2_W0_clk),
    .W0_data(mem_67_2_W0_data),
    .W0_en(mem_67_2_W0_en),
    .W0_mask(mem_67_2_W0_mask)
  );
  split_mem_0_ext mem_67_3 (
    .R0_addr(mem_67_3_R0_addr),
    .R0_clk(mem_67_3_R0_clk),
    .R0_data(mem_67_3_R0_data),
    .R0_en(mem_67_3_R0_en),
    .W0_addr(mem_67_3_W0_addr),
    .W0_clk(mem_67_3_W0_clk),
    .W0_data(mem_67_3_W0_data),
    .W0_en(mem_67_3_W0_en),
    .W0_mask(mem_67_3_W0_mask)
  );
  split_mem_0_ext mem_67_4 (
    .R0_addr(mem_67_4_R0_addr),
    .R0_clk(mem_67_4_R0_clk),
    .R0_data(mem_67_4_R0_data),
    .R0_en(mem_67_4_R0_en),
    .W0_addr(mem_67_4_W0_addr),
    .W0_clk(mem_67_4_W0_clk),
    .W0_data(mem_67_4_W0_data),
    .W0_en(mem_67_4_W0_en),
    .W0_mask(mem_67_4_W0_mask)
  );
  split_mem_0_ext mem_67_5 (
    .R0_addr(mem_67_5_R0_addr),
    .R0_clk(mem_67_5_R0_clk),
    .R0_data(mem_67_5_R0_data),
    .R0_en(mem_67_5_R0_en),
    .W0_addr(mem_67_5_W0_addr),
    .W0_clk(mem_67_5_W0_clk),
    .W0_data(mem_67_5_W0_data),
    .W0_en(mem_67_5_W0_en),
    .W0_mask(mem_67_5_W0_mask)
  );
  split_mem_0_ext mem_67_6 (
    .R0_addr(mem_67_6_R0_addr),
    .R0_clk(mem_67_6_R0_clk),
    .R0_data(mem_67_6_R0_data),
    .R0_en(mem_67_6_R0_en),
    .W0_addr(mem_67_6_W0_addr),
    .W0_clk(mem_67_6_W0_clk),
    .W0_data(mem_67_6_W0_data),
    .W0_en(mem_67_6_W0_en),
    .W0_mask(mem_67_6_W0_mask)
  );
  split_mem_0_ext mem_67_7 (
    .R0_addr(mem_67_7_R0_addr),
    .R0_clk(mem_67_7_R0_clk),
    .R0_data(mem_67_7_R0_data),
    .R0_en(mem_67_7_R0_en),
    .W0_addr(mem_67_7_W0_addr),
    .W0_clk(mem_67_7_W0_clk),
    .W0_data(mem_67_7_W0_data),
    .W0_en(mem_67_7_W0_en),
    .W0_mask(mem_67_7_W0_mask)
  );
  split_mem_0_ext mem_68_0 (
    .R0_addr(mem_68_0_R0_addr),
    .R0_clk(mem_68_0_R0_clk),
    .R0_data(mem_68_0_R0_data),
    .R0_en(mem_68_0_R0_en),
    .W0_addr(mem_68_0_W0_addr),
    .W0_clk(mem_68_0_W0_clk),
    .W0_data(mem_68_0_W0_data),
    .W0_en(mem_68_0_W0_en),
    .W0_mask(mem_68_0_W0_mask)
  );
  split_mem_0_ext mem_68_1 (
    .R0_addr(mem_68_1_R0_addr),
    .R0_clk(mem_68_1_R0_clk),
    .R0_data(mem_68_1_R0_data),
    .R0_en(mem_68_1_R0_en),
    .W0_addr(mem_68_1_W0_addr),
    .W0_clk(mem_68_1_W0_clk),
    .W0_data(mem_68_1_W0_data),
    .W0_en(mem_68_1_W0_en),
    .W0_mask(mem_68_1_W0_mask)
  );
  split_mem_0_ext mem_68_2 (
    .R0_addr(mem_68_2_R0_addr),
    .R0_clk(mem_68_2_R0_clk),
    .R0_data(mem_68_2_R0_data),
    .R0_en(mem_68_2_R0_en),
    .W0_addr(mem_68_2_W0_addr),
    .W0_clk(mem_68_2_W0_clk),
    .W0_data(mem_68_2_W0_data),
    .W0_en(mem_68_2_W0_en),
    .W0_mask(mem_68_2_W0_mask)
  );
  split_mem_0_ext mem_68_3 (
    .R0_addr(mem_68_3_R0_addr),
    .R0_clk(mem_68_3_R0_clk),
    .R0_data(mem_68_3_R0_data),
    .R0_en(mem_68_3_R0_en),
    .W0_addr(mem_68_3_W0_addr),
    .W0_clk(mem_68_3_W0_clk),
    .W0_data(mem_68_3_W0_data),
    .W0_en(mem_68_3_W0_en),
    .W0_mask(mem_68_3_W0_mask)
  );
  split_mem_0_ext mem_68_4 (
    .R0_addr(mem_68_4_R0_addr),
    .R0_clk(mem_68_4_R0_clk),
    .R0_data(mem_68_4_R0_data),
    .R0_en(mem_68_4_R0_en),
    .W0_addr(mem_68_4_W0_addr),
    .W0_clk(mem_68_4_W0_clk),
    .W0_data(mem_68_4_W0_data),
    .W0_en(mem_68_4_W0_en),
    .W0_mask(mem_68_4_W0_mask)
  );
  split_mem_0_ext mem_68_5 (
    .R0_addr(mem_68_5_R0_addr),
    .R0_clk(mem_68_5_R0_clk),
    .R0_data(mem_68_5_R0_data),
    .R0_en(mem_68_5_R0_en),
    .W0_addr(mem_68_5_W0_addr),
    .W0_clk(mem_68_5_W0_clk),
    .W0_data(mem_68_5_W0_data),
    .W0_en(mem_68_5_W0_en),
    .W0_mask(mem_68_5_W0_mask)
  );
  split_mem_0_ext mem_68_6 (
    .R0_addr(mem_68_6_R0_addr),
    .R0_clk(mem_68_6_R0_clk),
    .R0_data(mem_68_6_R0_data),
    .R0_en(mem_68_6_R0_en),
    .W0_addr(mem_68_6_W0_addr),
    .W0_clk(mem_68_6_W0_clk),
    .W0_data(mem_68_6_W0_data),
    .W0_en(mem_68_6_W0_en),
    .W0_mask(mem_68_6_W0_mask)
  );
  split_mem_0_ext mem_68_7 (
    .R0_addr(mem_68_7_R0_addr),
    .R0_clk(mem_68_7_R0_clk),
    .R0_data(mem_68_7_R0_data),
    .R0_en(mem_68_7_R0_en),
    .W0_addr(mem_68_7_W0_addr),
    .W0_clk(mem_68_7_W0_clk),
    .W0_data(mem_68_7_W0_data),
    .W0_en(mem_68_7_W0_en),
    .W0_mask(mem_68_7_W0_mask)
  );
  split_mem_0_ext mem_69_0 (
    .R0_addr(mem_69_0_R0_addr),
    .R0_clk(mem_69_0_R0_clk),
    .R0_data(mem_69_0_R0_data),
    .R0_en(mem_69_0_R0_en),
    .W0_addr(mem_69_0_W0_addr),
    .W0_clk(mem_69_0_W0_clk),
    .W0_data(mem_69_0_W0_data),
    .W0_en(mem_69_0_W0_en),
    .W0_mask(mem_69_0_W0_mask)
  );
  split_mem_0_ext mem_69_1 (
    .R0_addr(mem_69_1_R0_addr),
    .R0_clk(mem_69_1_R0_clk),
    .R0_data(mem_69_1_R0_data),
    .R0_en(mem_69_1_R0_en),
    .W0_addr(mem_69_1_W0_addr),
    .W0_clk(mem_69_1_W0_clk),
    .W0_data(mem_69_1_W0_data),
    .W0_en(mem_69_1_W0_en),
    .W0_mask(mem_69_1_W0_mask)
  );
  split_mem_0_ext mem_69_2 (
    .R0_addr(mem_69_2_R0_addr),
    .R0_clk(mem_69_2_R0_clk),
    .R0_data(mem_69_2_R0_data),
    .R0_en(mem_69_2_R0_en),
    .W0_addr(mem_69_2_W0_addr),
    .W0_clk(mem_69_2_W0_clk),
    .W0_data(mem_69_2_W0_data),
    .W0_en(mem_69_2_W0_en),
    .W0_mask(mem_69_2_W0_mask)
  );
  split_mem_0_ext mem_69_3 (
    .R0_addr(mem_69_3_R0_addr),
    .R0_clk(mem_69_3_R0_clk),
    .R0_data(mem_69_3_R0_data),
    .R0_en(mem_69_3_R0_en),
    .W0_addr(mem_69_3_W0_addr),
    .W0_clk(mem_69_3_W0_clk),
    .W0_data(mem_69_3_W0_data),
    .W0_en(mem_69_3_W0_en),
    .W0_mask(mem_69_3_W0_mask)
  );
  split_mem_0_ext mem_69_4 (
    .R0_addr(mem_69_4_R0_addr),
    .R0_clk(mem_69_4_R0_clk),
    .R0_data(mem_69_4_R0_data),
    .R0_en(mem_69_4_R0_en),
    .W0_addr(mem_69_4_W0_addr),
    .W0_clk(mem_69_4_W0_clk),
    .W0_data(mem_69_4_W0_data),
    .W0_en(mem_69_4_W0_en),
    .W0_mask(mem_69_4_W0_mask)
  );
  split_mem_0_ext mem_69_5 (
    .R0_addr(mem_69_5_R0_addr),
    .R0_clk(mem_69_5_R0_clk),
    .R0_data(mem_69_5_R0_data),
    .R0_en(mem_69_5_R0_en),
    .W0_addr(mem_69_5_W0_addr),
    .W0_clk(mem_69_5_W0_clk),
    .W0_data(mem_69_5_W0_data),
    .W0_en(mem_69_5_W0_en),
    .W0_mask(mem_69_5_W0_mask)
  );
  split_mem_0_ext mem_69_6 (
    .R0_addr(mem_69_6_R0_addr),
    .R0_clk(mem_69_6_R0_clk),
    .R0_data(mem_69_6_R0_data),
    .R0_en(mem_69_6_R0_en),
    .W0_addr(mem_69_6_W0_addr),
    .W0_clk(mem_69_6_W0_clk),
    .W0_data(mem_69_6_W0_data),
    .W0_en(mem_69_6_W0_en),
    .W0_mask(mem_69_6_W0_mask)
  );
  split_mem_0_ext mem_69_7 (
    .R0_addr(mem_69_7_R0_addr),
    .R0_clk(mem_69_7_R0_clk),
    .R0_data(mem_69_7_R0_data),
    .R0_en(mem_69_7_R0_en),
    .W0_addr(mem_69_7_W0_addr),
    .W0_clk(mem_69_7_W0_clk),
    .W0_data(mem_69_7_W0_data),
    .W0_en(mem_69_7_W0_en),
    .W0_mask(mem_69_7_W0_mask)
  );
  split_mem_0_ext mem_70_0 (
    .R0_addr(mem_70_0_R0_addr),
    .R0_clk(mem_70_0_R0_clk),
    .R0_data(mem_70_0_R0_data),
    .R0_en(mem_70_0_R0_en),
    .W0_addr(mem_70_0_W0_addr),
    .W0_clk(mem_70_0_W0_clk),
    .W0_data(mem_70_0_W0_data),
    .W0_en(mem_70_0_W0_en),
    .W0_mask(mem_70_0_W0_mask)
  );
  split_mem_0_ext mem_70_1 (
    .R0_addr(mem_70_1_R0_addr),
    .R0_clk(mem_70_1_R0_clk),
    .R0_data(mem_70_1_R0_data),
    .R0_en(mem_70_1_R0_en),
    .W0_addr(mem_70_1_W0_addr),
    .W0_clk(mem_70_1_W0_clk),
    .W0_data(mem_70_1_W0_data),
    .W0_en(mem_70_1_W0_en),
    .W0_mask(mem_70_1_W0_mask)
  );
  split_mem_0_ext mem_70_2 (
    .R0_addr(mem_70_2_R0_addr),
    .R0_clk(mem_70_2_R0_clk),
    .R0_data(mem_70_2_R0_data),
    .R0_en(mem_70_2_R0_en),
    .W0_addr(mem_70_2_W0_addr),
    .W0_clk(mem_70_2_W0_clk),
    .W0_data(mem_70_2_W0_data),
    .W0_en(mem_70_2_W0_en),
    .W0_mask(mem_70_2_W0_mask)
  );
  split_mem_0_ext mem_70_3 (
    .R0_addr(mem_70_3_R0_addr),
    .R0_clk(mem_70_3_R0_clk),
    .R0_data(mem_70_3_R0_data),
    .R0_en(mem_70_3_R0_en),
    .W0_addr(mem_70_3_W0_addr),
    .W0_clk(mem_70_3_W0_clk),
    .W0_data(mem_70_3_W0_data),
    .W0_en(mem_70_3_W0_en),
    .W0_mask(mem_70_3_W0_mask)
  );
  split_mem_0_ext mem_70_4 (
    .R0_addr(mem_70_4_R0_addr),
    .R0_clk(mem_70_4_R0_clk),
    .R0_data(mem_70_4_R0_data),
    .R0_en(mem_70_4_R0_en),
    .W0_addr(mem_70_4_W0_addr),
    .W0_clk(mem_70_4_W0_clk),
    .W0_data(mem_70_4_W0_data),
    .W0_en(mem_70_4_W0_en),
    .W0_mask(mem_70_4_W0_mask)
  );
  split_mem_0_ext mem_70_5 (
    .R0_addr(mem_70_5_R0_addr),
    .R0_clk(mem_70_5_R0_clk),
    .R0_data(mem_70_5_R0_data),
    .R0_en(mem_70_5_R0_en),
    .W0_addr(mem_70_5_W0_addr),
    .W0_clk(mem_70_5_W0_clk),
    .W0_data(mem_70_5_W0_data),
    .W0_en(mem_70_5_W0_en),
    .W0_mask(mem_70_5_W0_mask)
  );
  split_mem_0_ext mem_70_6 (
    .R0_addr(mem_70_6_R0_addr),
    .R0_clk(mem_70_6_R0_clk),
    .R0_data(mem_70_6_R0_data),
    .R0_en(mem_70_6_R0_en),
    .W0_addr(mem_70_6_W0_addr),
    .W0_clk(mem_70_6_W0_clk),
    .W0_data(mem_70_6_W0_data),
    .W0_en(mem_70_6_W0_en),
    .W0_mask(mem_70_6_W0_mask)
  );
  split_mem_0_ext mem_70_7 (
    .R0_addr(mem_70_7_R0_addr),
    .R0_clk(mem_70_7_R0_clk),
    .R0_data(mem_70_7_R0_data),
    .R0_en(mem_70_7_R0_en),
    .W0_addr(mem_70_7_W0_addr),
    .W0_clk(mem_70_7_W0_clk),
    .W0_data(mem_70_7_W0_data),
    .W0_en(mem_70_7_W0_en),
    .W0_mask(mem_70_7_W0_mask)
  );
  split_mem_0_ext mem_71_0 (
    .R0_addr(mem_71_0_R0_addr),
    .R0_clk(mem_71_0_R0_clk),
    .R0_data(mem_71_0_R0_data),
    .R0_en(mem_71_0_R0_en),
    .W0_addr(mem_71_0_W0_addr),
    .W0_clk(mem_71_0_W0_clk),
    .W0_data(mem_71_0_W0_data),
    .W0_en(mem_71_0_W0_en),
    .W0_mask(mem_71_0_W0_mask)
  );
  split_mem_0_ext mem_71_1 (
    .R0_addr(mem_71_1_R0_addr),
    .R0_clk(mem_71_1_R0_clk),
    .R0_data(mem_71_1_R0_data),
    .R0_en(mem_71_1_R0_en),
    .W0_addr(mem_71_1_W0_addr),
    .W0_clk(mem_71_1_W0_clk),
    .W0_data(mem_71_1_W0_data),
    .W0_en(mem_71_1_W0_en),
    .W0_mask(mem_71_1_W0_mask)
  );
  split_mem_0_ext mem_71_2 (
    .R0_addr(mem_71_2_R0_addr),
    .R0_clk(mem_71_2_R0_clk),
    .R0_data(mem_71_2_R0_data),
    .R0_en(mem_71_2_R0_en),
    .W0_addr(mem_71_2_W0_addr),
    .W0_clk(mem_71_2_W0_clk),
    .W0_data(mem_71_2_W0_data),
    .W0_en(mem_71_2_W0_en),
    .W0_mask(mem_71_2_W0_mask)
  );
  split_mem_0_ext mem_71_3 (
    .R0_addr(mem_71_3_R0_addr),
    .R0_clk(mem_71_3_R0_clk),
    .R0_data(mem_71_3_R0_data),
    .R0_en(mem_71_3_R0_en),
    .W0_addr(mem_71_3_W0_addr),
    .W0_clk(mem_71_3_W0_clk),
    .W0_data(mem_71_3_W0_data),
    .W0_en(mem_71_3_W0_en),
    .W0_mask(mem_71_3_W0_mask)
  );
  split_mem_0_ext mem_71_4 (
    .R0_addr(mem_71_4_R0_addr),
    .R0_clk(mem_71_4_R0_clk),
    .R0_data(mem_71_4_R0_data),
    .R0_en(mem_71_4_R0_en),
    .W0_addr(mem_71_4_W0_addr),
    .W0_clk(mem_71_4_W0_clk),
    .W0_data(mem_71_4_W0_data),
    .W0_en(mem_71_4_W0_en),
    .W0_mask(mem_71_4_W0_mask)
  );
  split_mem_0_ext mem_71_5 (
    .R0_addr(mem_71_5_R0_addr),
    .R0_clk(mem_71_5_R0_clk),
    .R0_data(mem_71_5_R0_data),
    .R0_en(mem_71_5_R0_en),
    .W0_addr(mem_71_5_W0_addr),
    .W0_clk(mem_71_5_W0_clk),
    .W0_data(mem_71_5_W0_data),
    .W0_en(mem_71_5_W0_en),
    .W0_mask(mem_71_5_W0_mask)
  );
  split_mem_0_ext mem_71_6 (
    .R0_addr(mem_71_6_R0_addr),
    .R0_clk(mem_71_6_R0_clk),
    .R0_data(mem_71_6_R0_data),
    .R0_en(mem_71_6_R0_en),
    .W0_addr(mem_71_6_W0_addr),
    .W0_clk(mem_71_6_W0_clk),
    .W0_data(mem_71_6_W0_data),
    .W0_en(mem_71_6_W0_en),
    .W0_mask(mem_71_6_W0_mask)
  );
  split_mem_0_ext mem_71_7 (
    .R0_addr(mem_71_7_R0_addr),
    .R0_clk(mem_71_7_R0_clk),
    .R0_data(mem_71_7_R0_data),
    .R0_en(mem_71_7_R0_en),
    .W0_addr(mem_71_7_W0_addr),
    .W0_clk(mem_71_7_W0_clk),
    .W0_data(mem_71_7_W0_data),
    .W0_en(mem_71_7_W0_en),
    .W0_mask(mem_71_7_W0_mask)
  );
  split_mem_0_ext mem_72_0 (
    .R0_addr(mem_72_0_R0_addr),
    .R0_clk(mem_72_0_R0_clk),
    .R0_data(mem_72_0_R0_data),
    .R0_en(mem_72_0_R0_en),
    .W0_addr(mem_72_0_W0_addr),
    .W0_clk(mem_72_0_W0_clk),
    .W0_data(mem_72_0_W0_data),
    .W0_en(mem_72_0_W0_en),
    .W0_mask(mem_72_0_W0_mask)
  );
  split_mem_0_ext mem_72_1 (
    .R0_addr(mem_72_1_R0_addr),
    .R0_clk(mem_72_1_R0_clk),
    .R0_data(mem_72_1_R0_data),
    .R0_en(mem_72_1_R0_en),
    .W0_addr(mem_72_1_W0_addr),
    .W0_clk(mem_72_1_W0_clk),
    .W0_data(mem_72_1_W0_data),
    .W0_en(mem_72_1_W0_en),
    .W0_mask(mem_72_1_W0_mask)
  );
  split_mem_0_ext mem_72_2 (
    .R0_addr(mem_72_2_R0_addr),
    .R0_clk(mem_72_2_R0_clk),
    .R0_data(mem_72_2_R0_data),
    .R0_en(mem_72_2_R0_en),
    .W0_addr(mem_72_2_W0_addr),
    .W0_clk(mem_72_2_W0_clk),
    .W0_data(mem_72_2_W0_data),
    .W0_en(mem_72_2_W0_en),
    .W0_mask(mem_72_2_W0_mask)
  );
  split_mem_0_ext mem_72_3 (
    .R0_addr(mem_72_3_R0_addr),
    .R0_clk(mem_72_3_R0_clk),
    .R0_data(mem_72_3_R0_data),
    .R0_en(mem_72_3_R0_en),
    .W0_addr(mem_72_3_W0_addr),
    .W0_clk(mem_72_3_W0_clk),
    .W0_data(mem_72_3_W0_data),
    .W0_en(mem_72_3_W0_en),
    .W0_mask(mem_72_3_W0_mask)
  );
  split_mem_0_ext mem_72_4 (
    .R0_addr(mem_72_4_R0_addr),
    .R0_clk(mem_72_4_R0_clk),
    .R0_data(mem_72_4_R0_data),
    .R0_en(mem_72_4_R0_en),
    .W0_addr(mem_72_4_W0_addr),
    .W0_clk(mem_72_4_W0_clk),
    .W0_data(mem_72_4_W0_data),
    .W0_en(mem_72_4_W0_en),
    .W0_mask(mem_72_4_W0_mask)
  );
  split_mem_0_ext mem_72_5 (
    .R0_addr(mem_72_5_R0_addr),
    .R0_clk(mem_72_5_R0_clk),
    .R0_data(mem_72_5_R0_data),
    .R0_en(mem_72_5_R0_en),
    .W0_addr(mem_72_5_W0_addr),
    .W0_clk(mem_72_5_W0_clk),
    .W0_data(mem_72_5_W0_data),
    .W0_en(mem_72_5_W0_en),
    .W0_mask(mem_72_5_W0_mask)
  );
  split_mem_0_ext mem_72_6 (
    .R0_addr(mem_72_6_R0_addr),
    .R0_clk(mem_72_6_R0_clk),
    .R0_data(mem_72_6_R0_data),
    .R0_en(mem_72_6_R0_en),
    .W0_addr(mem_72_6_W0_addr),
    .W0_clk(mem_72_6_W0_clk),
    .W0_data(mem_72_6_W0_data),
    .W0_en(mem_72_6_W0_en),
    .W0_mask(mem_72_6_W0_mask)
  );
  split_mem_0_ext mem_72_7 (
    .R0_addr(mem_72_7_R0_addr),
    .R0_clk(mem_72_7_R0_clk),
    .R0_data(mem_72_7_R0_data),
    .R0_en(mem_72_7_R0_en),
    .W0_addr(mem_72_7_W0_addr),
    .W0_clk(mem_72_7_W0_clk),
    .W0_data(mem_72_7_W0_data),
    .W0_en(mem_72_7_W0_en),
    .W0_mask(mem_72_7_W0_mask)
  );
  split_mem_0_ext mem_73_0 (
    .R0_addr(mem_73_0_R0_addr),
    .R0_clk(mem_73_0_R0_clk),
    .R0_data(mem_73_0_R0_data),
    .R0_en(mem_73_0_R0_en),
    .W0_addr(mem_73_0_W0_addr),
    .W0_clk(mem_73_0_W0_clk),
    .W0_data(mem_73_0_W0_data),
    .W0_en(mem_73_0_W0_en),
    .W0_mask(mem_73_0_W0_mask)
  );
  split_mem_0_ext mem_73_1 (
    .R0_addr(mem_73_1_R0_addr),
    .R0_clk(mem_73_1_R0_clk),
    .R0_data(mem_73_1_R0_data),
    .R0_en(mem_73_1_R0_en),
    .W0_addr(mem_73_1_W0_addr),
    .W0_clk(mem_73_1_W0_clk),
    .W0_data(mem_73_1_W0_data),
    .W0_en(mem_73_1_W0_en),
    .W0_mask(mem_73_1_W0_mask)
  );
  split_mem_0_ext mem_73_2 (
    .R0_addr(mem_73_2_R0_addr),
    .R0_clk(mem_73_2_R0_clk),
    .R0_data(mem_73_2_R0_data),
    .R0_en(mem_73_2_R0_en),
    .W0_addr(mem_73_2_W0_addr),
    .W0_clk(mem_73_2_W0_clk),
    .W0_data(mem_73_2_W0_data),
    .W0_en(mem_73_2_W0_en),
    .W0_mask(mem_73_2_W0_mask)
  );
  split_mem_0_ext mem_73_3 (
    .R0_addr(mem_73_3_R0_addr),
    .R0_clk(mem_73_3_R0_clk),
    .R0_data(mem_73_3_R0_data),
    .R0_en(mem_73_3_R0_en),
    .W0_addr(mem_73_3_W0_addr),
    .W0_clk(mem_73_3_W0_clk),
    .W0_data(mem_73_3_W0_data),
    .W0_en(mem_73_3_W0_en),
    .W0_mask(mem_73_3_W0_mask)
  );
  split_mem_0_ext mem_73_4 (
    .R0_addr(mem_73_4_R0_addr),
    .R0_clk(mem_73_4_R0_clk),
    .R0_data(mem_73_4_R0_data),
    .R0_en(mem_73_4_R0_en),
    .W0_addr(mem_73_4_W0_addr),
    .W0_clk(mem_73_4_W0_clk),
    .W0_data(mem_73_4_W0_data),
    .W0_en(mem_73_4_W0_en),
    .W0_mask(mem_73_4_W0_mask)
  );
  split_mem_0_ext mem_73_5 (
    .R0_addr(mem_73_5_R0_addr),
    .R0_clk(mem_73_5_R0_clk),
    .R0_data(mem_73_5_R0_data),
    .R0_en(mem_73_5_R0_en),
    .W0_addr(mem_73_5_W0_addr),
    .W0_clk(mem_73_5_W0_clk),
    .W0_data(mem_73_5_W0_data),
    .W0_en(mem_73_5_W0_en),
    .W0_mask(mem_73_5_W0_mask)
  );
  split_mem_0_ext mem_73_6 (
    .R0_addr(mem_73_6_R0_addr),
    .R0_clk(mem_73_6_R0_clk),
    .R0_data(mem_73_6_R0_data),
    .R0_en(mem_73_6_R0_en),
    .W0_addr(mem_73_6_W0_addr),
    .W0_clk(mem_73_6_W0_clk),
    .W0_data(mem_73_6_W0_data),
    .W0_en(mem_73_6_W0_en),
    .W0_mask(mem_73_6_W0_mask)
  );
  split_mem_0_ext mem_73_7 (
    .R0_addr(mem_73_7_R0_addr),
    .R0_clk(mem_73_7_R0_clk),
    .R0_data(mem_73_7_R0_data),
    .R0_en(mem_73_7_R0_en),
    .W0_addr(mem_73_7_W0_addr),
    .W0_clk(mem_73_7_W0_clk),
    .W0_data(mem_73_7_W0_data),
    .W0_en(mem_73_7_W0_en),
    .W0_mask(mem_73_7_W0_mask)
  );
  split_mem_0_ext mem_74_0 (
    .R0_addr(mem_74_0_R0_addr),
    .R0_clk(mem_74_0_R0_clk),
    .R0_data(mem_74_0_R0_data),
    .R0_en(mem_74_0_R0_en),
    .W0_addr(mem_74_0_W0_addr),
    .W0_clk(mem_74_0_W0_clk),
    .W0_data(mem_74_0_W0_data),
    .W0_en(mem_74_0_W0_en),
    .W0_mask(mem_74_0_W0_mask)
  );
  split_mem_0_ext mem_74_1 (
    .R0_addr(mem_74_1_R0_addr),
    .R0_clk(mem_74_1_R0_clk),
    .R0_data(mem_74_1_R0_data),
    .R0_en(mem_74_1_R0_en),
    .W0_addr(mem_74_1_W0_addr),
    .W0_clk(mem_74_1_W0_clk),
    .W0_data(mem_74_1_W0_data),
    .W0_en(mem_74_1_W0_en),
    .W0_mask(mem_74_1_W0_mask)
  );
  split_mem_0_ext mem_74_2 (
    .R0_addr(mem_74_2_R0_addr),
    .R0_clk(mem_74_2_R0_clk),
    .R0_data(mem_74_2_R0_data),
    .R0_en(mem_74_2_R0_en),
    .W0_addr(mem_74_2_W0_addr),
    .W0_clk(mem_74_2_W0_clk),
    .W0_data(mem_74_2_W0_data),
    .W0_en(mem_74_2_W0_en),
    .W0_mask(mem_74_2_W0_mask)
  );
  split_mem_0_ext mem_74_3 (
    .R0_addr(mem_74_3_R0_addr),
    .R0_clk(mem_74_3_R0_clk),
    .R0_data(mem_74_3_R0_data),
    .R0_en(mem_74_3_R0_en),
    .W0_addr(mem_74_3_W0_addr),
    .W0_clk(mem_74_3_W0_clk),
    .W0_data(mem_74_3_W0_data),
    .W0_en(mem_74_3_W0_en),
    .W0_mask(mem_74_3_W0_mask)
  );
  split_mem_0_ext mem_74_4 (
    .R0_addr(mem_74_4_R0_addr),
    .R0_clk(mem_74_4_R0_clk),
    .R0_data(mem_74_4_R0_data),
    .R0_en(mem_74_4_R0_en),
    .W0_addr(mem_74_4_W0_addr),
    .W0_clk(mem_74_4_W0_clk),
    .W0_data(mem_74_4_W0_data),
    .W0_en(mem_74_4_W0_en),
    .W0_mask(mem_74_4_W0_mask)
  );
  split_mem_0_ext mem_74_5 (
    .R0_addr(mem_74_5_R0_addr),
    .R0_clk(mem_74_5_R0_clk),
    .R0_data(mem_74_5_R0_data),
    .R0_en(mem_74_5_R0_en),
    .W0_addr(mem_74_5_W0_addr),
    .W0_clk(mem_74_5_W0_clk),
    .W0_data(mem_74_5_W0_data),
    .W0_en(mem_74_5_W0_en),
    .W0_mask(mem_74_5_W0_mask)
  );
  split_mem_0_ext mem_74_6 (
    .R0_addr(mem_74_6_R0_addr),
    .R0_clk(mem_74_6_R0_clk),
    .R0_data(mem_74_6_R0_data),
    .R0_en(mem_74_6_R0_en),
    .W0_addr(mem_74_6_W0_addr),
    .W0_clk(mem_74_6_W0_clk),
    .W0_data(mem_74_6_W0_data),
    .W0_en(mem_74_6_W0_en),
    .W0_mask(mem_74_6_W0_mask)
  );
  split_mem_0_ext mem_74_7 (
    .R0_addr(mem_74_7_R0_addr),
    .R0_clk(mem_74_7_R0_clk),
    .R0_data(mem_74_7_R0_data),
    .R0_en(mem_74_7_R0_en),
    .W0_addr(mem_74_7_W0_addr),
    .W0_clk(mem_74_7_W0_clk),
    .W0_data(mem_74_7_W0_data),
    .W0_en(mem_74_7_W0_en),
    .W0_mask(mem_74_7_W0_mask)
  );
  split_mem_0_ext mem_75_0 (
    .R0_addr(mem_75_0_R0_addr),
    .R0_clk(mem_75_0_R0_clk),
    .R0_data(mem_75_0_R0_data),
    .R0_en(mem_75_0_R0_en),
    .W0_addr(mem_75_0_W0_addr),
    .W0_clk(mem_75_0_W0_clk),
    .W0_data(mem_75_0_W0_data),
    .W0_en(mem_75_0_W0_en),
    .W0_mask(mem_75_0_W0_mask)
  );
  split_mem_0_ext mem_75_1 (
    .R0_addr(mem_75_1_R0_addr),
    .R0_clk(mem_75_1_R0_clk),
    .R0_data(mem_75_1_R0_data),
    .R0_en(mem_75_1_R0_en),
    .W0_addr(mem_75_1_W0_addr),
    .W0_clk(mem_75_1_W0_clk),
    .W0_data(mem_75_1_W0_data),
    .W0_en(mem_75_1_W0_en),
    .W0_mask(mem_75_1_W0_mask)
  );
  split_mem_0_ext mem_75_2 (
    .R0_addr(mem_75_2_R0_addr),
    .R0_clk(mem_75_2_R0_clk),
    .R0_data(mem_75_2_R0_data),
    .R0_en(mem_75_2_R0_en),
    .W0_addr(mem_75_2_W0_addr),
    .W0_clk(mem_75_2_W0_clk),
    .W0_data(mem_75_2_W0_data),
    .W0_en(mem_75_2_W0_en),
    .W0_mask(mem_75_2_W0_mask)
  );
  split_mem_0_ext mem_75_3 (
    .R0_addr(mem_75_3_R0_addr),
    .R0_clk(mem_75_3_R0_clk),
    .R0_data(mem_75_3_R0_data),
    .R0_en(mem_75_3_R0_en),
    .W0_addr(mem_75_3_W0_addr),
    .W0_clk(mem_75_3_W0_clk),
    .W0_data(mem_75_3_W0_data),
    .W0_en(mem_75_3_W0_en),
    .W0_mask(mem_75_3_W0_mask)
  );
  split_mem_0_ext mem_75_4 (
    .R0_addr(mem_75_4_R0_addr),
    .R0_clk(mem_75_4_R0_clk),
    .R0_data(mem_75_4_R0_data),
    .R0_en(mem_75_4_R0_en),
    .W0_addr(mem_75_4_W0_addr),
    .W0_clk(mem_75_4_W0_clk),
    .W0_data(mem_75_4_W0_data),
    .W0_en(mem_75_4_W0_en),
    .W0_mask(mem_75_4_W0_mask)
  );
  split_mem_0_ext mem_75_5 (
    .R0_addr(mem_75_5_R0_addr),
    .R0_clk(mem_75_5_R0_clk),
    .R0_data(mem_75_5_R0_data),
    .R0_en(mem_75_5_R0_en),
    .W0_addr(mem_75_5_W0_addr),
    .W0_clk(mem_75_5_W0_clk),
    .W0_data(mem_75_5_W0_data),
    .W0_en(mem_75_5_W0_en),
    .W0_mask(mem_75_5_W0_mask)
  );
  split_mem_0_ext mem_75_6 (
    .R0_addr(mem_75_6_R0_addr),
    .R0_clk(mem_75_6_R0_clk),
    .R0_data(mem_75_6_R0_data),
    .R0_en(mem_75_6_R0_en),
    .W0_addr(mem_75_6_W0_addr),
    .W0_clk(mem_75_6_W0_clk),
    .W0_data(mem_75_6_W0_data),
    .W0_en(mem_75_6_W0_en),
    .W0_mask(mem_75_6_W0_mask)
  );
  split_mem_0_ext mem_75_7 (
    .R0_addr(mem_75_7_R0_addr),
    .R0_clk(mem_75_7_R0_clk),
    .R0_data(mem_75_7_R0_data),
    .R0_en(mem_75_7_R0_en),
    .W0_addr(mem_75_7_W0_addr),
    .W0_clk(mem_75_7_W0_clk),
    .W0_data(mem_75_7_W0_data),
    .W0_en(mem_75_7_W0_en),
    .W0_mask(mem_75_7_W0_mask)
  );
  split_mem_0_ext mem_76_0 (
    .R0_addr(mem_76_0_R0_addr),
    .R0_clk(mem_76_0_R0_clk),
    .R0_data(mem_76_0_R0_data),
    .R0_en(mem_76_0_R0_en),
    .W0_addr(mem_76_0_W0_addr),
    .W0_clk(mem_76_0_W0_clk),
    .W0_data(mem_76_0_W0_data),
    .W0_en(mem_76_0_W0_en),
    .W0_mask(mem_76_0_W0_mask)
  );
  split_mem_0_ext mem_76_1 (
    .R0_addr(mem_76_1_R0_addr),
    .R0_clk(mem_76_1_R0_clk),
    .R0_data(mem_76_1_R0_data),
    .R0_en(mem_76_1_R0_en),
    .W0_addr(mem_76_1_W0_addr),
    .W0_clk(mem_76_1_W0_clk),
    .W0_data(mem_76_1_W0_data),
    .W0_en(mem_76_1_W0_en),
    .W0_mask(mem_76_1_W0_mask)
  );
  split_mem_0_ext mem_76_2 (
    .R0_addr(mem_76_2_R0_addr),
    .R0_clk(mem_76_2_R0_clk),
    .R0_data(mem_76_2_R0_data),
    .R0_en(mem_76_2_R0_en),
    .W0_addr(mem_76_2_W0_addr),
    .W0_clk(mem_76_2_W0_clk),
    .W0_data(mem_76_2_W0_data),
    .W0_en(mem_76_2_W0_en),
    .W0_mask(mem_76_2_W0_mask)
  );
  split_mem_0_ext mem_76_3 (
    .R0_addr(mem_76_3_R0_addr),
    .R0_clk(mem_76_3_R0_clk),
    .R0_data(mem_76_3_R0_data),
    .R0_en(mem_76_3_R0_en),
    .W0_addr(mem_76_3_W0_addr),
    .W0_clk(mem_76_3_W0_clk),
    .W0_data(mem_76_3_W0_data),
    .W0_en(mem_76_3_W0_en),
    .W0_mask(mem_76_3_W0_mask)
  );
  split_mem_0_ext mem_76_4 (
    .R0_addr(mem_76_4_R0_addr),
    .R0_clk(mem_76_4_R0_clk),
    .R0_data(mem_76_4_R0_data),
    .R0_en(mem_76_4_R0_en),
    .W0_addr(mem_76_4_W0_addr),
    .W0_clk(mem_76_4_W0_clk),
    .W0_data(mem_76_4_W0_data),
    .W0_en(mem_76_4_W0_en),
    .W0_mask(mem_76_4_W0_mask)
  );
  split_mem_0_ext mem_76_5 (
    .R0_addr(mem_76_5_R0_addr),
    .R0_clk(mem_76_5_R0_clk),
    .R0_data(mem_76_5_R0_data),
    .R0_en(mem_76_5_R0_en),
    .W0_addr(mem_76_5_W0_addr),
    .W0_clk(mem_76_5_W0_clk),
    .W0_data(mem_76_5_W0_data),
    .W0_en(mem_76_5_W0_en),
    .W0_mask(mem_76_5_W0_mask)
  );
  split_mem_0_ext mem_76_6 (
    .R0_addr(mem_76_6_R0_addr),
    .R0_clk(mem_76_6_R0_clk),
    .R0_data(mem_76_6_R0_data),
    .R0_en(mem_76_6_R0_en),
    .W0_addr(mem_76_6_W0_addr),
    .W0_clk(mem_76_6_W0_clk),
    .W0_data(mem_76_6_W0_data),
    .W0_en(mem_76_6_W0_en),
    .W0_mask(mem_76_6_W0_mask)
  );
  split_mem_0_ext mem_76_7 (
    .R0_addr(mem_76_7_R0_addr),
    .R0_clk(mem_76_7_R0_clk),
    .R0_data(mem_76_7_R0_data),
    .R0_en(mem_76_7_R0_en),
    .W0_addr(mem_76_7_W0_addr),
    .W0_clk(mem_76_7_W0_clk),
    .W0_data(mem_76_7_W0_data),
    .W0_en(mem_76_7_W0_en),
    .W0_mask(mem_76_7_W0_mask)
  );
  split_mem_0_ext mem_77_0 (
    .R0_addr(mem_77_0_R0_addr),
    .R0_clk(mem_77_0_R0_clk),
    .R0_data(mem_77_0_R0_data),
    .R0_en(mem_77_0_R0_en),
    .W0_addr(mem_77_0_W0_addr),
    .W0_clk(mem_77_0_W0_clk),
    .W0_data(mem_77_0_W0_data),
    .W0_en(mem_77_0_W0_en),
    .W0_mask(mem_77_0_W0_mask)
  );
  split_mem_0_ext mem_77_1 (
    .R0_addr(mem_77_1_R0_addr),
    .R0_clk(mem_77_1_R0_clk),
    .R0_data(mem_77_1_R0_data),
    .R0_en(mem_77_1_R0_en),
    .W0_addr(mem_77_1_W0_addr),
    .W0_clk(mem_77_1_W0_clk),
    .W0_data(mem_77_1_W0_data),
    .W0_en(mem_77_1_W0_en),
    .W0_mask(mem_77_1_W0_mask)
  );
  split_mem_0_ext mem_77_2 (
    .R0_addr(mem_77_2_R0_addr),
    .R0_clk(mem_77_2_R0_clk),
    .R0_data(mem_77_2_R0_data),
    .R0_en(mem_77_2_R0_en),
    .W0_addr(mem_77_2_W0_addr),
    .W0_clk(mem_77_2_W0_clk),
    .W0_data(mem_77_2_W0_data),
    .W0_en(mem_77_2_W0_en),
    .W0_mask(mem_77_2_W0_mask)
  );
  split_mem_0_ext mem_77_3 (
    .R0_addr(mem_77_3_R0_addr),
    .R0_clk(mem_77_3_R0_clk),
    .R0_data(mem_77_3_R0_data),
    .R0_en(mem_77_3_R0_en),
    .W0_addr(mem_77_3_W0_addr),
    .W0_clk(mem_77_3_W0_clk),
    .W0_data(mem_77_3_W0_data),
    .W0_en(mem_77_3_W0_en),
    .W0_mask(mem_77_3_W0_mask)
  );
  split_mem_0_ext mem_77_4 (
    .R0_addr(mem_77_4_R0_addr),
    .R0_clk(mem_77_4_R0_clk),
    .R0_data(mem_77_4_R0_data),
    .R0_en(mem_77_4_R0_en),
    .W0_addr(mem_77_4_W0_addr),
    .W0_clk(mem_77_4_W0_clk),
    .W0_data(mem_77_4_W0_data),
    .W0_en(mem_77_4_W0_en),
    .W0_mask(mem_77_4_W0_mask)
  );
  split_mem_0_ext mem_77_5 (
    .R0_addr(mem_77_5_R0_addr),
    .R0_clk(mem_77_5_R0_clk),
    .R0_data(mem_77_5_R0_data),
    .R0_en(mem_77_5_R0_en),
    .W0_addr(mem_77_5_W0_addr),
    .W0_clk(mem_77_5_W0_clk),
    .W0_data(mem_77_5_W0_data),
    .W0_en(mem_77_5_W0_en),
    .W0_mask(mem_77_5_W0_mask)
  );
  split_mem_0_ext mem_77_6 (
    .R0_addr(mem_77_6_R0_addr),
    .R0_clk(mem_77_6_R0_clk),
    .R0_data(mem_77_6_R0_data),
    .R0_en(mem_77_6_R0_en),
    .W0_addr(mem_77_6_W0_addr),
    .W0_clk(mem_77_6_W0_clk),
    .W0_data(mem_77_6_W0_data),
    .W0_en(mem_77_6_W0_en),
    .W0_mask(mem_77_6_W0_mask)
  );
  split_mem_0_ext mem_77_7 (
    .R0_addr(mem_77_7_R0_addr),
    .R0_clk(mem_77_7_R0_clk),
    .R0_data(mem_77_7_R0_data),
    .R0_en(mem_77_7_R0_en),
    .W0_addr(mem_77_7_W0_addr),
    .W0_clk(mem_77_7_W0_clk),
    .W0_data(mem_77_7_W0_data),
    .W0_en(mem_77_7_W0_en),
    .W0_mask(mem_77_7_W0_mask)
  );
  split_mem_0_ext mem_78_0 (
    .R0_addr(mem_78_0_R0_addr),
    .R0_clk(mem_78_0_R0_clk),
    .R0_data(mem_78_0_R0_data),
    .R0_en(mem_78_0_R0_en),
    .W0_addr(mem_78_0_W0_addr),
    .W0_clk(mem_78_0_W0_clk),
    .W0_data(mem_78_0_W0_data),
    .W0_en(mem_78_0_W0_en),
    .W0_mask(mem_78_0_W0_mask)
  );
  split_mem_0_ext mem_78_1 (
    .R0_addr(mem_78_1_R0_addr),
    .R0_clk(mem_78_1_R0_clk),
    .R0_data(mem_78_1_R0_data),
    .R0_en(mem_78_1_R0_en),
    .W0_addr(mem_78_1_W0_addr),
    .W0_clk(mem_78_1_W0_clk),
    .W0_data(mem_78_1_W0_data),
    .W0_en(mem_78_1_W0_en),
    .W0_mask(mem_78_1_W0_mask)
  );
  split_mem_0_ext mem_78_2 (
    .R0_addr(mem_78_2_R0_addr),
    .R0_clk(mem_78_2_R0_clk),
    .R0_data(mem_78_2_R0_data),
    .R0_en(mem_78_2_R0_en),
    .W0_addr(mem_78_2_W0_addr),
    .W0_clk(mem_78_2_W0_clk),
    .W0_data(mem_78_2_W0_data),
    .W0_en(mem_78_2_W0_en),
    .W0_mask(mem_78_2_W0_mask)
  );
  split_mem_0_ext mem_78_3 (
    .R0_addr(mem_78_3_R0_addr),
    .R0_clk(mem_78_3_R0_clk),
    .R0_data(mem_78_3_R0_data),
    .R0_en(mem_78_3_R0_en),
    .W0_addr(mem_78_3_W0_addr),
    .W0_clk(mem_78_3_W0_clk),
    .W0_data(mem_78_3_W0_data),
    .W0_en(mem_78_3_W0_en),
    .W0_mask(mem_78_3_W0_mask)
  );
  split_mem_0_ext mem_78_4 (
    .R0_addr(mem_78_4_R0_addr),
    .R0_clk(mem_78_4_R0_clk),
    .R0_data(mem_78_4_R0_data),
    .R0_en(mem_78_4_R0_en),
    .W0_addr(mem_78_4_W0_addr),
    .W0_clk(mem_78_4_W0_clk),
    .W0_data(mem_78_4_W0_data),
    .W0_en(mem_78_4_W0_en),
    .W0_mask(mem_78_4_W0_mask)
  );
  split_mem_0_ext mem_78_5 (
    .R0_addr(mem_78_5_R0_addr),
    .R0_clk(mem_78_5_R0_clk),
    .R0_data(mem_78_5_R0_data),
    .R0_en(mem_78_5_R0_en),
    .W0_addr(mem_78_5_W0_addr),
    .W0_clk(mem_78_5_W0_clk),
    .W0_data(mem_78_5_W0_data),
    .W0_en(mem_78_5_W0_en),
    .W0_mask(mem_78_5_W0_mask)
  );
  split_mem_0_ext mem_78_6 (
    .R0_addr(mem_78_6_R0_addr),
    .R0_clk(mem_78_6_R0_clk),
    .R0_data(mem_78_6_R0_data),
    .R0_en(mem_78_6_R0_en),
    .W0_addr(mem_78_6_W0_addr),
    .W0_clk(mem_78_6_W0_clk),
    .W0_data(mem_78_6_W0_data),
    .W0_en(mem_78_6_W0_en),
    .W0_mask(mem_78_6_W0_mask)
  );
  split_mem_0_ext mem_78_7 (
    .R0_addr(mem_78_7_R0_addr),
    .R0_clk(mem_78_7_R0_clk),
    .R0_data(mem_78_7_R0_data),
    .R0_en(mem_78_7_R0_en),
    .W0_addr(mem_78_7_W0_addr),
    .W0_clk(mem_78_7_W0_clk),
    .W0_data(mem_78_7_W0_data),
    .W0_en(mem_78_7_W0_en),
    .W0_mask(mem_78_7_W0_mask)
  );
  split_mem_0_ext mem_79_0 (
    .R0_addr(mem_79_0_R0_addr),
    .R0_clk(mem_79_0_R0_clk),
    .R0_data(mem_79_0_R0_data),
    .R0_en(mem_79_0_R0_en),
    .W0_addr(mem_79_0_W0_addr),
    .W0_clk(mem_79_0_W0_clk),
    .W0_data(mem_79_0_W0_data),
    .W0_en(mem_79_0_W0_en),
    .W0_mask(mem_79_0_W0_mask)
  );
  split_mem_0_ext mem_79_1 (
    .R0_addr(mem_79_1_R0_addr),
    .R0_clk(mem_79_1_R0_clk),
    .R0_data(mem_79_1_R0_data),
    .R0_en(mem_79_1_R0_en),
    .W0_addr(mem_79_1_W0_addr),
    .W0_clk(mem_79_1_W0_clk),
    .W0_data(mem_79_1_W0_data),
    .W0_en(mem_79_1_W0_en),
    .W0_mask(mem_79_1_W0_mask)
  );
  split_mem_0_ext mem_79_2 (
    .R0_addr(mem_79_2_R0_addr),
    .R0_clk(mem_79_2_R0_clk),
    .R0_data(mem_79_2_R0_data),
    .R0_en(mem_79_2_R0_en),
    .W0_addr(mem_79_2_W0_addr),
    .W0_clk(mem_79_2_W0_clk),
    .W0_data(mem_79_2_W0_data),
    .W0_en(mem_79_2_W0_en),
    .W0_mask(mem_79_2_W0_mask)
  );
  split_mem_0_ext mem_79_3 (
    .R0_addr(mem_79_3_R0_addr),
    .R0_clk(mem_79_3_R0_clk),
    .R0_data(mem_79_3_R0_data),
    .R0_en(mem_79_3_R0_en),
    .W0_addr(mem_79_3_W0_addr),
    .W0_clk(mem_79_3_W0_clk),
    .W0_data(mem_79_3_W0_data),
    .W0_en(mem_79_3_W0_en),
    .W0_mask(mem_79_3_W0_mask)
  );
  split_mem_0_ext mem_79_4 (
    .R0_addr(mem_79_4_R0_addr),
    .R0_clk(mem_79_4_R0_clk),
    .R0_data(mem_79_4_R0_data),
    .R0_en(mem_79_4_R0_en),
    .W0_addr(mem_79_4_W0_addr),
    .W0_clk(mem_79_4_W0_clk),
    .W0_data(mem_79_4_W0_data),
    .W0_en(mem_79_4_W0_en),
    .W0_mask(mem_79_4_W0_mask)
  );
  split_mem_0_ext mem_79_5 (
    .R0_addr(mem_79_5_R0_addr),
    .R0_clk(mem_79_5_R0_clk),
    .R0_data(mem_79_5_R0_data),
    .R0_en(mem_79_5_R0_en),
    .W0_addr(mem_79_5_W0_addr),
    .W0_clk(mem_79_5_W0_clk),
    .W0_data(mem_79_5_W0_data),
    .W0_en(mem_79_5_W0_en),
    .W0_mask(mem_79_5_W0_mask)
  );
  split_mem_0_ext mem_79_6 (
    .R0_addr(mem_79_6_R0_addr),
    .R0_clk(mem_79_6_R0_clk),
    .R0_data(mem_79_6_R0_data),
    .R0_en(mem_79_6_R0_en),
    .W0_addr(mem_79_6_W0_addr),
    .W0_clk(mem_79_6_W0_clk),
    .W0_data(mem_79_6_W0_data),
    .W0_en(mem_79_6_W0_en),
    .W0_mask(mem_79_6_W0_mask)
  );
  split_mem_0_ext mem_79_7 (
    .R0_addr(mem_79_7_R0_addr),
    .R0_clk(mem_79_7_R0_clk),
    .R0_data(mem_79_7_R0_data),
    .R0_en(mem_79_7_R0_en),
    .W0_addr(mem_79_7_W0_addr),
    .W0_clk(mem_79_7_W0_clk),
    .W0_data(mem_79_7_W0_data),
    .W0_en(mem_79_7_W0_en),
    .W0_mask(mem_79_7_W0_mask)
  );
  split_mem_0_ext mem_80_0 (
    .R0_addr(mem_80_0_R0_addr),
    .R0_clk(mem_80_0_R0_clk),
    .R0_data(mem_80_0_R0_data),
    .R0_en(mem_80_0_R0_en),
    .W0_addr(mem_80_0_W0_addr),
    .W0_clk(mem_80_0_W0_clk),
    .W0_data(mem_80_0_W0_data),
    .W0_en(mem_80_0_W0_en),
    .W0_mask(mem_80_0_W0_mask)
  );
  split_mem_0_ext mem_80_1 (
    .R0_addr(mem_80_1_R0_addr),
    .R0_clk(mem_80_1_R0_clk),
    .R0_data(mem_80_1_R0_data),
    .R0_en(mem_80_1_R0_en),
    .W0_addr(mem_80_1_W0_addr),
    .W0_clk(mem_80_1_W0_clk),
    .W0_data(mem_80_1_W0_data),
    .W0_en(mem_80_1_W0_en),
    .W0_mask(mem_80_1_W0_mask)
  );
  split_mem_0_ext mem_80_2 (
    .R0_addr(mem_80_2_R0_addr),
    .R0_clk(mem_80_2_R0_clk),
    .R0_data(mem_80_2_R0_data),
    .R0_en(mem_80_2_R0_en),
    .W0_addr(mem_80_2_W0_addr),
    .W0_clk(mem_80_2_W0_clk),
    .W0_data(mem_80_2_W0_data),
    .W0_en(mem_80_2_W0_en),
    .W0_mask(mem_80_2_W0_mask)
  );
  split_mem_0_ext mem_80_3 (
    .R0_addr(mem_80_3_R0_addr),
    .R0_clk(mem_80_3_R0_clk),
    .R0_data(mem_80_3_R0_data),
    .R0_en(mem_80_3_R0_en),
    .W0_addr(mem_80_3_W0_addr),
    .W0_clk(mem_80_3_W0_clk),
    .W0_data(mem_80_3_W0_data),
    .W0_en(mem_80_3_W0_en),
    .W0_mask(mem_80_3_W0_mask)
  );
  split_mem_0_ext mem_80_4 (
    .R0_addr(mem_80_4_R0_addr),
    .R0_clk(mem_80_4_R0_clk),
    .R0_data(mem_80_4_R0_data),
    .R0_en(mem_80_4_R0_en),
    .W0_addr(mem_80_4_W0_addr),
    .W0_clk(mem_80_4_W0_clk),
    .W0_data(mem_80_4_W0_data),
    .W0_en(mem_80_4_W0_en),
    .W0_mask(mem_80_4_W0_mask)
  );
  split_mem_0_ext mem_80_5 (
    .R0_addr(mem_80_5_R0_addr),
    .R0_clk(mem_80_5_R0_clk),
    .R0_data(mem_80_5_R0_data),
    .R0_en(mem_80_5_R0_en),
    .W0_addr(mem_80_5_W0_addr),
    .W0_clk(mem_80_5_W0_clk),
    .W0_data(mem_80_5_W0_data),
    .W0_en(mem_80_5_W0_en),
    .W0_mask(mem_80_5_W0_mask)
  );
  split_mem_0_ext mem_80_6 (
    .R0_addr(mem_80_6_R0_addr),
    .R0_clk(mem_80_6_R0_clk),
    .R0_data(mem_80_6_R0_data),
    .R0_en(mem_80_6_R0_en),
    .W0_addr(mem_80_6_W0_addr),
    .W0_clk(mem_80_6_W0_clk),
    .W0_data(mem_80_6_W0_data),
    .W0_en(mem_80_6_W0_en),
    .W0_mask(mem_80_6_W0_mask)
  );
  split_mem_0_ext mem_80_7 (
    .R0_addr(mem_80_7_R0_addr),
    .R0_clk(mem_80_7_R0_clk),
    .R0_data(mem_80_7_R0_data),
    .R0_en(mem_80_7_R0_en),
    .W0_addr(mem_80_7_W0_addr),
    .W0_clk(mem_80_7_W0_clk),
    .W0_data(mem_80_7_W0_data),
    .W0_en(mem_80_7_W0_en),
    .W0_mask(mem_80_7_W0_mask)
  );
  split_mem_0_ext mem_81_0 (
    .R0_addr(mem_81_0_R0_addr),
    .R0_clk(mem_81_0_R0_clk),
    .R0_data(mem_81_0_R0_data),
    .R0_en(mem_81_0_R0_en),
    .W0_addr(mem_81_0_W0_addr),
    .W0_clk(mem_81_0_W0_clk),
    .W0_data(mem_81_0_W0_data),
    .W0_en(mem_81_0_W0_en),
    .W0_mask(mem_81_0_W0_mask)
  );
  split_mem_0_ext mem_81_1 (
    .R0_addr(mem_81_1_R0_addr),
    .R0_clk(mem_81_1_R0_clk),
    .R0_data(mem_81_1_R0_data),
    .R0_en(mem_81_1_R0_en),
    .W0_addr(mem_81_1_W0_addr),
    .W0_clk(mem_81_1_W0_clk),
    .W0_data(mem_81_1_W0_data),
    .W0_en(mem_81_1_W0_en),
    .W0_mask(mem_81_1_W0_mask)
  );
  split_mem_0_ext mem_81_2 (
    .R0_addr(mem_81_2_R0_addr),
    .R0_clk(mem_81_2_R0_clk),
    .R0_data(mem_81_2_R0_data),
    .R0_en(mem_81_2_R0_en),
    .W0_addr(mem_81_2_W0_addr),
    .W0_clk(mem_81_2_W0_clk),
    .W0_data(mem_81_2_W0_data),
    .W0_en(mem_81_2_W0_en),
    .W0_mask(mem_81_2_W0_mask)
  );
  split_mem_0_ext mem_81_3 (
    .R0_addr(mem_81_3_R0_addr),
    .R0_clk(mem_81_3_R0_clk),
    .R0_data(mem_81_3_R0_data),
    .R0_en(mem_81_3_R0_en),
    .W0_addr(mem_81_3_W0_addr),
    .W0_clk(mem_81_3_W0_clk),
    .W0_data(mem_81_3_W0_data),
    .W0_en(mem_81_3_W0_en),
    .W0_mask(mem_81_3_W0_mask)
  );
  split_mem_0_ext mem_81_4 (
    .R0_addr(mem_81_4_R0_addr),
    .R0_clk(mem_81_4_R0_clk),
    .R0_data(mem_81_4_R0_data),
    .R0_en(mem_81_4_R0_en),
    .W0_addr(mem_81_4_W0_addr),
    .W0_clk(mem_81_4_W0_clk),
    .W0_data(mem_81_4_W0_data),
    .W0_en(mem_81_4_W0_en),
    .W0_mask(mem_81_4_W0_mask)
  );
  split_mem_0_ext mem_81_5 (
    .R0_addr(mem_81_5_R0_addr),
    .R0_clk(mem_81_5_R0_clk),
    .R0_data(mem_81_5_R0_data),
    .R0_en(mem_81_5_R0_en),
    .W0_addr(mem_81_5_W0_addr),
    .W0_clk(mem_81_5_W0_clk),
    .W0_data(mem_81_5_W0_data),
    .W0_en(mem_81_5_W0_en),
    .W0_mask(mem_81_5_W0_mask)
  );
  split_mem_0_ext mem_81_6 (
    .R0_addr(mem_81_6_R0_addr),
    .R0_clk(mem_81_6_R0_clk),
    .R0_data(mem_81_6_R0_data),
    .R0_en(mem_81_6_R0_en),
    .W0_addr(mem_81_6_W0_addr),
    .W0_clk(mem_81_6_W0_clk),
    .W0_data(mem_81_6_W0_data),
    .W0_en(mem_81_6_W0_en),
    .W0_mask(mem_81_6_W0_mask)
  );
  split_mem_0_ext mem_81_7 (
    .R0_addr(mem_81_7_R0_addr),
    .R0_clk(mem_81_7_R0_clk),
    .R0_data(mem_81_7_R0_data),
    .R0_en(mem_81_7_R0_en),
    .W0_addr(mem_81_7_W0_addr),
    .W0_clk(mem_81_7_W0_clk),
    .W0_data(mem_81_7_W0_data),
    .W0_en(mem_81_7_W0_en),
    .W0_mask(mem_81_7_W0_mask)
  );
  split_mem_0_ext mem_82_0 (
    .R0_addr(mem_82_0_R0_addr),
    .R0_clk(mem_82_0_R0_clk),
    .R0_data(mem_82_0_R0_data),
    .R0_en(mem_82_0_R0_en),
    .W0_addr(mem_82_0_W0_addr),
    .W0_clk(mem_82_0_W0_clk),
    .W0_data(mem_82_0_W0_data),
    .W0_en(mem_82_0_W0_en),
    .W0_mask(mem_82_0_W0_mask)
  );
  split_mem_0_ext mem_82_1 (
    .R0_addr(mem_82_1_R0_addr),
    .R0_clk(mem_82_1_R0_clk),
    .R0_data(mem_82_1_R0_data),
    .R0_en(mem_82_1_R0_en),
    .W0_addr(mem_82_1_W0_addr),
    .W0_clk(mem_82_1_W0_clk),
    .W0_data(mem_82_1_W0_data),
    .W0_en(mem_82_1_W0_en),
    .W0_mask(mem_82_1_W0_mask)
  );
  split_mem_0_ext mem_82_2 (
    .R0_addr(mem_82_2_R0_addr),
    .R0_clk(mem_82_2_R0_clk),
    .R0_data(mem_82_2_R0_data),
    .R0_en(mem_82_2_R0_en),
    .W0_addr(mem_82_2_W0_addr),
    .W0_clk(mem_82_2_W0_clk),
    .W0_data(mem_82_2_W0_data),
    .W0_en(mem_82_2_W0_en),
    .W0_mask(mem_82_2_W0_mask)
  );
  split_mem_0_ext mem_82_3 (
    .R0_addr(mem_82_3_R0_addr),
    .R0_clk(mem_82_3_R0_clk),
    .R0_data(mem_82_3_R0_data),
    .R0_en(mem_82_3_R0_en),
    .W0_addr(mem_82_3_W0_addr),
    .W0_clk(mem_82_3_W0_clk),
    .W0_data(mem_82_3_W0_data),
    .W0_en(mem_82_3_W0_en),
    .W0_mask(mem_82_3_W0_mask)
  );
  split_mem_0_ext mem_82_4 (
    .R0_addr(mem_82_4_R0_addr),
    .R0_clk(mem_82_4_R0_clk),
    .R0_data(mem_82_4_R0_data),
    .R0_en(mem_82_4_R0_en),
    .W0_addr(mem_82_4_W0_addr),
    .W0_clk(mem_82_4_W0_clk),
    .W0_data(mem_82_4_W0_data),
    .W0_en(mem_82_4_W0_en),
    .W0_mask(mem_82_4_W0_mask)
  );
  split_mem_0_ext mem_82_5 (
    .R0_addr(mem_82_5_R0_addr),
    .R0_clk(mem_82_5_R0_clk),
    .R0_data(mem_82_5_R0_data),
    .R0_en(mem_82_5_R0_en),
    .W0_addr(mem_82_5_W0_addr),
    .W0_clk(mem_82_5_W0_clk),
    .W0_data(mem_82_5_W0_data),
    .W0_en(mem_82_5_W0_en),
    .W0_mask(mem_82_5_W0_mask)
  );
  split_mem_0_ext mem_82_6 (
    .R0_addr(mem_82_6_R0_addr),
    .R0_clk(mem_82_6_R0_clk),
    .R0_data(mem_82_6_R0_data),
    .R0_en(mem_82_6_R0_en),
    .W0_addr(mem_82_6_W0_addr),
    .W0_clk(mem_82_6_W0_clk),
    .W0_data(mem_82_6_W0_data),
    .W0_en(mem_82_6_W0_en),
    .W0_mask(mem_82_6_W0_mask)
  );
  split_mem_0_ext mem_82_7 (
    .R0_addr(mem_82_7_R0_addr),
    .R0_clk(mem_82_7_R0_clk),
    .R0_data(mem_82_7_R0_data),
    .R0_en(mem_82_7_R0_en),
    .W0_addr(mem_82_7_W0_addr),
    .W0_clk(mem_82_7_W0_clk),
    .W0_data(mem_82_7_W0_data),
    .W0_en(mem_82_7_W0_en),
    .W0_mask(mem_82_7_W0_mask)
  );
  split_mem_0_ext mem_83_0 (
    .R0_addr(mem_83_0_R0_addr),
    .R0_clk(mem_83_0_R0_clk),
    .R0_data(mem_83_0_R0_data),
    .R0_en(mem_83_0_R0_en),
    .W0_addr(mem_83_0_W0_addr),
    .W0_clk(mem_83_0_W0_clk),
    .W0_data(mem_83_0_W0_data),
    .W0_en(mem_83_0_W0_en),
    .W0_mask(mem_83_0_W0_mask)
  );
  split_mem_0_ext mem_83_1 (
    .R0_addr(mem_83_1_R0_addr),
    .R0_clk(mem_83_1_R0_clk),
    .R0_data(mem_83_1_R0_data),
    .R0_en(mem_83_1_R0_en),
    .W0_addr(mem_83_1_W0_addr),
    .W0_clk(mem_83_1_W0_clk),
    .W0_data(mem_83_1_W0_data),
    .W0_en(mem_83_1_W0_en),
    .W0_mask(mem_83_1_W0_mask)
  );
  split_mem_0_ext mem_83_2 (
    .R0_addr(mem_83_2_R0_addr),
    .R0_clk(mem_83_2_R0_clk),
    .R0_data(mem_83_2_R0_data),
    .R0_en(mem_83_2_R0_en),
    .W0_addr(mem_83_2_W0_addr),
    .W0_clk(mem_83_2_W0_clk),
    .W0_data(mem_83_2_W0_data),
    .W0_en(mem_83_2_W0_en),
    .W0_mask(mem_83_2_W0_mask)
  );
  split_mem_0_ext mem_83_3 (
    .R0_addr(mem_83_3_R0_addr),
    .R0_clk(mem_83_3_R0_clk),
    .R0_data(mem_83_3_R0_data),
    .R0_en(mem_83_3_R0_en),
    .W0_addr(mem_83_3_W0_addr),
    .W0_clk(mem_83_3_W0_clk),
    .W0_data(mem_83_3_W0_data),
    .W0_en(mem_83_3_W0_en),
    .W0_mask(mem_83_3_W0_mask)
  );
  split_mem_0_ext mem_83_4 (
    .R0_addr(mem_83_4_R0_addr),
    .R0_clk(mem_83_4_R0_clk),
    .R0_data(mem_83_4_R0_data),
    .R0_en(mem_83_4_R0_en),
    .W0_addr(mem_83_4_W0_addr),
    .W0_clk(mem_83_4_W0_clk),
    .W0_data(mem_83_4_W0_data),
    .W0_en(mem_83_4_W0_en),
    .W0_mask(mem_83_4_W0_mask)
  );
  split_mem_0_ext mem_83_5 (
    .R0_addr(mem_83_5_R0_addr),
    .R0_clk(mem_83_5_R0_clk),
    .R0_data(mem_83_5_R0_data),
    .R0_en(mem_83_5_R0_en),
    .W0_addr(mem_83_5_W0_addr),
    .W0_clk(mem_83_5_W0_clk),
    .W0_data(mem_83_5_W0_data),
    .W0_en(mem_83_5_W0_en),
    .W0_mask(mem_83_5_W0_mask)
  );
  split_mem_0_ext mem_83_6 (
    .R0_addr(mem_83_6_R0_addr),
    .R0_clk(mem_83_6_R0_clk),
    .R0_data(mem_83_6_R0_data),
    .R0_en(mem_83_6_R0_en),
    .W0_addr(mem_83_6_W0_addr),
    .W0_clk(mem_83_6_W0_clk),
    .W0_data(mem_83_6_W0_data),
    .W0_en(mem_83_6_W0_en),
    .W0_mask(mem_83_6_W0_mask)
  );
  split_mem_0_ext mem_83_7 (
    .R0_addr(mem_83_7_R0_addr),
    .R0_clk(mem_83_7_R0_clk),
    .R0_data(mem_83_7_R0_data),
    .R0_en(mem_83_7_R0_en),
    .W0_addr(mem_83_7_W0_addr),
    .W0_clk(mem_83_7_W0_clk),
    .W0_data(mem_83_7_W0_data),
    .W0_en(mem_83_7_W0_en),
    .W0_mask(mem_83_7_W0_mask)
  );
  split_mem_0_ext mem_84_0 (
    .R0_addr(mem_84_0_R0_addr),
    .R0_clk(mem_84_0_R0_clk),
    .R0_data(mem_84_0_R0_data),
    .R0_en(mem_84_0_R0_en),
    .W0_addr(mem_84_0_W0_addr),
    .W0_clk(mem_84_0_W0_clk),
    .W0_data(mem_84_0_W0_data),
    .W0_en(mem_84_0_W0_en),
    .W0_mask(mem_84_0_W0_mask)
  );
  split_mem_0_ext mem_84_1 (
    .R0_addr(mem_84_1_R0_addr),
    .R0_clk(mem_84_1_R0_clk),
    .R0_data(mem_84_1_R0_data),
    .R0_en(mem_84_1_R0_en),
    .W0_addr(mem_84_1_W0_addr),
    .W0_clk(mem_84_1_W0_clk),
    .W0_data(mem_84_1_W0_data),
    .W0_en(mem_84_1_W0_en),
    .W0_mask(mem_84_1_W0_mask)
  );
  split_mem_0_ext mem_84_2 (
    .R0_addr(mem_84_2_R0_addr),
    .R0_clk(mem_84_2_R0_clk),
    .R0_data(mem_84_2_R0_data),
    .R0_en(mem_84_2_R0_en),
    .W0_addr(mem_84_2_W0_addr),
    .W0_clk(mem_84_2_W0_clk),
    .W0_data(mem_84_2_W0_data),
    .W0_en(mem_84_2_W0_en),
    .W0_mask(mem_84_2_W0_mask)
  );
  split_mem_0_ext mem_84_3 (
    .R0_addr(mem_84_3_R0_addr),
    .R0_clk(mem_84_3_R0_clk),
    .R0_data(mem_84_3_R0_data),
    .R0_en(mem_84_3_R0_en),
    .W0_addr(mem_84_3_W0_addr),
    .W0_clk(mem_84_3_W0_clk),
    .W0_data(mem_84_3_W0_data),
    .W0_en(mem_84_3_W0_en),
    .W0_mask(mem_84_3_W0_mask)
  );
  split_mem_0_ext mem_84_4 (
    .R0_addr(mem_84_4_R0_addr),
    .R0_clk(mem_84_4_R0_clk),
    .R0_data(mem_84_4_R0_data),
    .R0_en(mem_84_4_R0_en),
    .W0_addr(mem_84_4_W0_addr),
    .W0_clk(mem_84_4_W0_clk),
    .W0_data(mem_84_4_W0_data),
    .W0_en(mem_84_4_W0_en),
    .W0_mask(mem_84_4_W0_mask)
  );
  split_mem_0_ext mem_84_5 (
    .R0_addr(mem_84_5_R0_addr),
    .R0_clk(mem_84_5_R0_clk),
    .R0_data(mem_84_5_R0_data),
    .R0_en(mem_84_5_R0_en),
    .W0_addr(mem_84_5_W0_addr),
    .W0_clk(mem_84_5_W0_clk),
    .W0_data(mem_84_5_W0_data),
    .W0_en(mem_84_5_W0_en),
    .W0_mask(mem_84_5_W0_mask)
  );
  split_mem_0_ext mem_84_6 (
    .R0_addr(mem_84_6_R0_addr),
    .R0_clk(mem_84_6_R0_clk),
    .R0_data(mem_84_6_R0_data),
    .R0_en(mem_84_6_R0_en),
    .W0_addr(mem_84_6_W0_addr),
    .W0_clk(mem_84_6_W0_clk),
    .W0_data(mem_84_6_W0_data),
    .W0_en(mem_84_6_W0_en),
    .W0_mask(mem_84_6_W0_mask)
  );
  split_mem_0_ext mem_84_7 (
    .R0_addr(mem_84_7_R0_addr),
    .R0_clk(mem_84_7_R0_clk),
    .R0_data(mem_84_7_R0_data),
    .R0_en(mem_84_7_R0_en),
    .W0_addr(mem_84_7_W0_addr),
    .W0_clk(mem_84_7_W0_clk),
    .W0_data(mem_84_7_W0_data),
    .W0_en(mem_84_7_W0_en),
    .W0_mask(mem_84_7_W0_mask)
  );
  split_mem_0_ext mem_85_0 (
    .R0_addr(mem_85_0_R0_addr),
    .R0_clk(mem_85_0_R0_clk),
    .R0_data(mem_85_0_R0_data),
    .R0_en(mem_85_0_R0_en),
    .W0_addr(mem_85_0_W0_addr),
    .W0_clk(mem_85_0_W0_clk),
    .W0_data(mem_85_0_W0_data),
    .W0_en(mem_85_0_W0_en),
    .W0_mask(mem_85_0_W0_mask)
  );
  split_mem_0_ext mem_85_1 (
    .R0_addr(mem_85_1_R0_addr),
    .R0_clk(mem_85_1_R0_clk),
    .R0_data(mem_85_1_R0_data),
    .R0_en(mem_85_1_R0_en),
    .W0_addr(mem_85_1_W0_addr),
    .W0_clk(mem_85_1_W0_clk),
    .W0_data(mem_85_1_W0_data),
    .W0_en(mem_85_1_W0_en),
    .W0_mask(mem_85_1_W0_mask)
  );
  split_mem_0_ext mem_85_2 (
    .R0_addr(mem_85_2_R0_addr),
    .R0_clk(mem_85_2_R0_clk),
    .R0_data(mem_85_2_R0_data),
    .R0_en(mem_85_2_R0_en),
    .W0_addr(mem_85_2_W0_addr),
    .W0_clk(mem_85_2_W0_clk),
    .W0_data(mem_85_2_W0_data),
    .W0_en(mem_85_2_W0_en),
    .W0_mask(mem_85_2_W0_mask)
  );
  split_mem_0_ext mem_85_3 (
    .R0_addr(mem_85_3_R0_addr),
    .R0_clk(mem_85_3_R0_clk),
    .R0_data(mem_85_3_R0_data),
    .R0_en(mem_85_3_R0_en),
    .W0_addr(mem_85_3_W0_addr),
    .W0_clk(mem_85_3_W0_clk),
    .W0_data(mem_85_3_W0_data),
    .W0_en(mem_85_3_W0_en),
    .W0_mask(mem_85_3_W0_mask)
  );
  split_mem_0_ext mem_85_4 (
    .R0_addr(mem_85_4_R0_addr),
    .R0_clk(mem_85_4_R0_clk),
    .R0_data(mem_85_4_R0_data),
    .R0_en(mem_85_4_R0_en),
    .W0_addr(mem_85_4_W0_addr),
    .W0_clk(mem_85_4_W0_clk),
    .W0_data(mem_85_4_W0_data),
    .W0_en(mem_85_4_W0_en),
    .W0_mask(mem_85_4_W0_mask)
  );
  split_mem_0_ext mem_85_5 (
    .R0_addr(mem_85_5_R0_addr),
    .R0_clk(mem_85_5_R0_clk),
    .R0_data(mem_85_5_R0_data),
    .R0_en(mem_85_5_R0_en),
    .W0_addr(mem_85_5_W0_addr),
    .W0_clk(mem_85_5_W0_clk),
    .W0_data(mem_85_5_W0_data),
    .W0_en(mem_85_5_W0_en),
    .W0_mask(mem_85_5_W0_mask)
  );
  split_mem_0_ext mem_85_6 (
    .R0_addr(mem_85_6_R0_addr),
    .R0_clk(mem_85_6_R0_clk),
    .R0_data(mem_85_6_R0_data),
    .R0_en(mem_85_6_R0_en),
    .W0_addr(mem_85_6_W0_addr),
    .W0_clk(mem_85_6_W0_clk),
    .W0_data(mem_85_6_W0_data),
    .W0_en(mem_85_6_W0_en),
    .W0_mask(mem_85_6_W0_mask)
  );
  split_mem_0_ext mem_85_7 (
    .R0_addr(mem_85_7_R0_addr),
    .R0_clk(mem_85_7_R0_clk),
    .R0_data(mem_85_7_R0_data),
    .R0_en(mem_85_7_R0_en),
    .W0_addr(mem_85_7_W0_addr),
    .W0_clk(mem_85_7_W0_clk),
    .W0_data(mem_85_7_W0_data),
    .W0_en(mem_85_7_W0_en),
    .W0_mask(mem_85_7_W0_mask)
  );
  split_mem_0_ext mem_86_0 (
    .R0_addr(mem_86_0_R0_addr),
    .R0_clk(mem_86_0_R0_clk),
    .R0_data(mem_86_0_R0_data),
    .R0_en(mem_86_0_R0_en),
    .W0_addr(mem_86_0_W0_addr),
    .W0_clk(mem_86_0_W0_clk),
    .W0_data(mem_86_0_W0_data),
    .W0_en(mem_86_0_W0_en),
    .W0_mask(mem_86_0_W0_mask)
  );
  split_mem_0_ext mem_86_1 (
    .R0_addr(mem_86_1_R0_addr),
    .R0_clk(mem_86_1_R0_clk),
    .R0_data(mem_86_1_R0_data),
    .R0_en(mem_86_1_R0_en),
    .W0_addr(mem_86_1_W0_addr),
    .W0_clk(mem_86_1_W0_clk),
    .W0_data(mem_86_1_W0_data),
    .W0_en(mem_86_1_W0_en),
    .W0_mask(mem_86_1_W0_mask)
  );
  split_mem_0_ext mem_86_2 (
    .R0_addr(mem_86_2_R0_addr),
    .R0_clk(mem_86_2_R0_clk),
    .R0_data(mem_86_2_R0_data),
    .R0_en(mem_86_2_R0_en),
    .W0_addr(mem_86_2_W0_addr),
    .W0_clk(mem_86_2_W0_clk),
    .W0_data(mem_86_2_W0_data),
    .W0_en(mem_86_2_W0_en),
    .W0_mask(mem_86_2_W0_mask)
  );
  split_mem_0_ext mem_86_3 (
    .R0_addr(mem_86_3_R0_addr),
    .R0_clk(mem_86_3_R0_clk),
    .R0_data(mem_86_3_R0_data),
    .R0_en(mem_86_3_R0_en),
    .W0_addr(mem_86_3_W0_addr),
    .W0_clk(mem_86_3_W0_clk),
    .W0_data(mem_86_3_W0_data),
    .W0_en(mem_86_3_W0_en),
    .W0_mask(mem_86_3_W0_mask)
  );
  split_mem_0_ext mem_86_4 (
    .R0_addr(mem_86_4_R0_addr),
    .R0_clk(mem_86_4_R0_clk),
    .R0_data(mem_86_4_R0_data),
    .R0_en(mem_86_4_R0_en),
    .W0_addr(mem_86_4_W0_addr),
    .W0_clk(mem_86_4_W0_clk),
    .W0_data(mem_86_4_W0_data),
    .W0_en(mem_86_4_W0_en),
    .W0_mask(mem_86_4_W0_mask)
  );
  split_mem_0_ext mem_86_5 (
    .R0_addr(mem_86_5_R0_addr),
    .R0_clk(mem_86_5_R0_clk),
    .R0_data(mem_86_5_R0_data),
    .R0_en(mem_86_5_R0_en),
    .W0_addr(mem_86_5_W0_addr),
    .W0_clk(mem_86_5_W0_clk),
    .W0_data(mem_86_5_W0_data),
    .W0_en(mem_86_5_W0_en),
    .W0_mask(mem_86_5_W0_mask)
  );
  split_mem_0_ext mem_86_6 (
    .R0_addr(mem_86_6_R0_addr),
    .R0_clk(mem_86_6_R0_clk),
    .R0_data(mem_86_6_R0_data),
    .R0_en(mem_86_6_R0_en),
    .W0_addr(mem_86_6_W0_addr),
    .W0_clk(mem_86_6_W0_clk),
    .W0_data(mem_86_6_W0_data),
    .W0_en(mem_86_6_W0_en),
    .W0_mask(mem_86_6_W0_mask)
  );
  split_mem_0_ext mem_86_7 (
    .R0_addr(mem_86_7_R0_addr),
    .R0_clk(mem_86_7_R0_clk),
    .R0_data(mem_86_7_R0_data),
    .R0_en(mem_86_7_R0_en),
    .W0_addr(mem_86_7_W0_addr),
    .W0_clk(mem_86_7_W0_clk),
    .W0_data(mem_86_7_W0_data),
    .W0_en(mem_86_7_W0_en),
    .W0_mask(mem_86_7_W0_mask)
  );
  split_mem_0_ext mem_87_0 (
    .R0_addr(mem_87_0_R0_addr),
    .R0_clk(mem_87_0_R0_clk),
    .R0_data(mem_87_0_R0_data),
    .R0_en(mem_87_0_R0_en),
    .W0_addr(mem_87_0_W0_addr),
    .W0_clk(mem_87_0_W0_clk),
    .W0_data(mem_87_0_W0_data),
    .W0_en(mem_87_0_W0_en),
    .W0_mask(mem_87_0_W0_mask)
  );
  split_mem_0_ext mem_87_1 (
    .R0_addr(mem_87_1_R0_addr),
    .R0_clk(mem_87_1_R0_clk),
    .R0_data(mem_87_1_R0_data),
    .R0_en(mem_87_1_R0_en),
    .W0_addr(mem_87_1_W0_addr),
    .W0_clk(mem_87_1_W0_clk),
    .W0_data(mem_87_1_W0_data),
    .W0_en(mem_87_1_W0_en),
    .W0_mask(mem_87_1_W0_mask)
  );
  split_mem_0_ext mem_87_2 (
    .R0_addr(mem_87_2_R0_addr),
    .R0_clk(mem_87_2_R0_clk),
    .R0_data(mem_87_2_R0_data),
    .R0_en(mem_87_2_R0_en),
    .W0_addr(mem_87_2_W0_addr),
    .W0_clk(mem_87_2_W0_clk),
    .W0_data(mem_87_2_W0_data),
    .W0_en(mem_87_2_W0_en),
    .W0_mask(mem_87_2_W0_mask)
  );
  split_mem_0_ext mem_87_3 (
    .R0_addr(mem_87_3_R0_addr),
    .R0_clk(mem_87_3_R0_clk),
    .R0_data(mem_87_3_R0_data),
    .R0_en(mem_87_3_R0_en),
    .W0_addr(mem_87_3_W0_addr),
    .W0_clk(mem_87_3_W0_clk),
    .W0_data(mem_87_3_W0_data),
    .W0_en(mem_87_3_W0_en),
    .W0_mask(mem_87_3_W0_mask)
  );
  split_mem_0_ext mem_87_4 (
    .R0_addr(mem_87_4_R0_addr),
    .R0_clk(mem_87_4_R0_clk),
    .R0_data(mem_87_4_R0_data),
    .R0_en(mem_87_4_R0_en),
    .W0_addr(mem_87_4_W0_addr),
    .W0_clk(mem_87_4_W0_clk),
    .W0_data(mem_87_4_W0_data),
    .W0_en(mem_87_4_W0_en),
    .W0_mask(mem_87_4_W0_mask)
  );
  split_mem_0_ext mem_87_5 (
    .R0_addr(mem_87_5_R0_addr),
    .R0_clk(mem_87_5_R0_clk),
    .R0_data(mem_87_5_R0_data),
    .R0_en(mem_87_5_R0_en),
    .W0_addr(mem_87_5_W0_addr),
    .W0_clk(mem_87_5_W0_clk),
    .W0_data(mem_87_5_W0_data),
    .W0_en(mem_87_5_W0_en),
    .W0_mask(mem_87_5_W0_mask)
  );
  split_mem_0_ext mem_87_6 (
    .R0_addr(mem_87_6_R0_addr),
    .R0_clk(mem_87_6_R0_clk),
    .R0_data(mem_87_6_R0_data),
    .R0_en(mem_87_6_R0_en),
    .W0_addr(mem_87_6_W0_addr),
    .W0_clk(mem_87_6_W0_clk),
    .W0_data(mem_87_6_W0_data),
    .W0_en(mem_87_6_W0_en),
    .W0_mask(mem_87_6_W0_mask)
  );
  split_mem_0_ext mem_87_7 (
    .R0_addr(mem_87_7_R0_addr),
    .R0_clk(mem_87_7_R0_clk),
    .R0_data(mem_87_7_R0_data),
    .R0_en(mem_87_7_R0_en),
    .W0_addr(mem_87_7_W0_addr),
    .W0_clk(mem_87_7_W0_clk),
    .W0_data(mem_87_7_W0_data),
    .W0_en(mem_87_7_W0_en),
    .W0_mask(mem_87_7_W0_mask)
  );
  split_mem_0_ext mem_88_0 (
    .R0_addr(mem_88_0_R0_addr),
    .R0_clk(mem_88_0_R0_clk),
    .R0_data(mem_88_0_R0_data),
    .R0_en(mem_88_0_R0_en),
    .W0_addr(mem_88_0_W0_addr),
    .W0_clk(mem_88_0_W0_clk),
    .W0_data(mem_88_0_W0_data),
    .W0_en(mem_88_0_W0_en),
    .W0_mask(mem_88_0_W0_mask)
  );
  split_mem_0_ext mem_88_1 (
    .R0_addr(mem_88_1_R0_addr),
    .R0_clk(mem_88_1_R0_clk),
    .R0_data(mem_88_1_R0_data),
    .R0_en(mem_88_1_R0_en),
    .W0_addr(mem_88_1_W0_addr),
    .W0_clk(mem_88_1_W0_clk),
    .W0_data(mem_88_1_W0_data),
    .W0_en(mem_88_1_W0_en),
    .W0_mask(mem_88_1_W0_mask)
  );
  split_mem_0_ext mem_88_2 (
    .R0_addr(mem_88_2_R0_addr),
    .R0_clk(mem_88_2_R0_clk),
    .R0_data(mem_88_2_R0_data),
    .R0_en(mem_88_2_R0_en),
    .W0_addr(mem_88_2_W0_addr),
    .W0_clk(mem_88_2_W0_clk),
    .W0_data(mem_88_2_W0_data),
    .W0_en(mem_88_2_W0_en),
    .W0_mask(mem_88_2_W0_mask)
  );
  split_mem_0_ext mem_88_3 (
    .R0_addr(mem_88_3_R0_addr),
    .R0_clk(mem_88_3_R0_clk),
    .R0_data(mem_88_3_R0_data),
    .R0_en(mem_88_3_R0_en),
    .W0_addr(mem_88_3_W0_addr),
    .W0_clk(mem_88_3_W0_clk),
    .W0_data(mem_88_3_W0_data),
    .W0_en(mem_88_3_W0_en),
    .W0_mask(mem_88_3_W0_mask)
  );
  split_mem_0_ext mem_88_4 (
    .R0_addr(mem_88_4_R0_addr),
    .R0_clk(mem_88_4_R0_clk),
    .R0_data(mem_88_4_R0_data),
    .R0_en(mem_88_4_R0_en),
    .W0_addr(mem_88_4_W0_addr),
    .W0_clk(mem_88_4_W0_clk),
    .W0_data(mem_88_4_W0_data),
    .W0_en(mem_88_4_W0_en),
    .W0_mask(mem_88_4_W0_mask)
  );
  split_mem_0_ext mem_88_5 (
    .R0_addr(mem_88_5_R0_addr),
    .R0_clk(mem_88_5_R0_clk),
    .R0_data(mem_88_5_R0_data),
    .R0_en(mem_88_5_R0_en),
    .W0_addr(mem_88_5_W0_addr),
    .W0_clk(mem_88_5_W0_clk),
    .W0_data(mem_88_5_W0_data),
    .W0_en(mem_88_5_W0_en),
    .W0_mask(mem_88_5_W0_mask)
  );
  split_mem_0_ext mem_88_6 (
    .R0_addr(mem_88_6_R0_addr),
    .R0_clk(mem_88_6_R0_clk),
    .R0_data(mem_88_6_R0_data),
    .R0_en(mem_88_6_R0_en),
    .W0_addr(mem_88_6_W0_addr),
    .W0_clk(mem_88_6_W0_clk),
    .W0_data(mem_88_6_W0_data),
    .W0_en(mem_88_6_W0_en),
    .W0_mask(mem_88_6_W0_mask)
  );
  split_mem_0_ext mem_88_7 (
    .R0_addr(mem_88_7_R0_addr),
    .R0_clk(mem_88_7_R0_clk),
    .R0_data(mem_88_7_R0_data),
    .R0_en(mem_88_7_R0_en),
    .W0_addr(mem_88_7_W0_addr),
    .W0_clk(mem_88_7_W0_clk),
    .W0_data(mem_88_7_W0_data),
    .W0_en(mem_88_7_W0_en),
    .W0_mask(mem_88_7_W0_mask)
  );
  split_mem_0_ext mem_89_0 (
    .R0_addr(mem_89_0_R0_addr),
    .R0_clk(mem_89_0_R0_clk),
    .R0_data(mem_89_0_R0_data),
    .R0_en(mem_89_0_R0_en),
    .W0_addr(mem_89_0_W0_addr),
    .W0_clk(mem_89_0_W0_clk),
    .W0_data(mem_89_0_W0_data),
    .W0_en(mem_89_0_W0_en),
    .W0_mask(mem_89_0_W0_mask)
  );
  split_mem_0_ext mem_89_1 (
    .R0_addr(mem_89_1_R0_addr),
    .R0_clk(mem_89_1_R0_clk),
    .R0_data(mem_89_1_R0_data),
    .R0_en(mem_89_1_R0_en),
    .W0_addr(mem_89_1_W0_addr),
    .W0_clk(mem_89_1_W0_clk),
    .W0_data(mem_89_1_W0_data),
    .W0_en(mem_89_1_W0_en),
    .W0_mask(mem_89_1_W0_mask)
  );
  split_mem_0_ext mem_89_2 (
    .R0_addr(mem_89_2_R0_addr),
    .R0_clk(mem_89_2_R0_clk),
    .R0_data(mem_89_2_R0_data),
    .R0_en(mem_89_2_R0_en),
    .W0_addr(mem_89_2_W0_addr),
    .W0_clk(mem_89_2_W0_clk),
    .W0_data(mem_89_2_W0_data),
    .W0_en(mem_89_2_W0_en),
    .W0_mask(mem_89_2_W0_mask)
  );
  split_mem_0_ext mem_89_3 (
    .R0_addr(mem_89_3_R0_addr),
    .R0_clk(mem_89_3_R0_clk),
    .R0_data(mem_89_3_R0_data),
    .R0_en(mem_89_3_R0_en),
    .W0_addr(mem_89_3_W0_addr),
    .W0_clk(mem_89_3_W0_clk),
    .W0_data(mem_89_3_W0_data),
    .W0_en(mem_89_3_W0_en),
    .W0_mask(mem_89_3_W0_mask)
  );
  split_mem_0_ext mem_89_4 (
    .R0_addr(mem_89_4_R0_addr),
    .R0_clk(mem_89_4_R0_clk),
    .R0_data(mem_89_4_R0_data),
    .R0_en(mem_89_4_R0_en),
    .W0_addr(mem_89_4_W0_addr),
    .W0_clk(mem_89_4_W0_clk),
    .W0_data(mem_89_4_W0_data),
    .W0_en(mem_89_4_W0_en),
    .W0_mask(mem_89_4_W0_mask)
  );
  split_mem_0_ext mem_89_5 (
    .R0_addr(mem_89_5_R0_addr),
    .R0_clk(mem_89_5_R0_clk),
    .R0_data(mem_89_5_R0_data),
    .R0_en(mem_89_5_R0_en),
    .W0_addr(mem_89_5_W0_addr),
    .W0_clk(mem_89_5_W0_clk),
    .W0_data(mem_89_5_W0_data),
    .W0_en(mem_89_5_W0_en),
    .W0_mask(mem_89_5_W0_mask)
  );
  split_mem_0_ext mem_89_6 (
    .R0_addr(mem_89_6_R0_addr),
    .R0_clk(mem_89_6_R0_clk),
    .R0_data(mem_89_6_R0_data),
    .R0_en(mem_89_6_R0_en),
    .W0_addr(mem_89_6_W0_addr),
    .W0_clk(mem_89_6_W0_clk),
    .W0_data(mem_89_6_W0_data),
    .W0_en(mem_89_6_W0_en),
    .W0_mask(mem_89_6_W0_mask)
  );
  split_mem_0_ext mem_89_7 (
    .R0_addr(mem_89_7_R0_addr),
    .R0_clk(mem_89_7_R0_clk),
    .R0_data(mem_89_7_R0_data),
    .R0_en(mem_89_7_R0_en),
    .W0_addr(mem_89_7_W0_addr),
    .W0_clk(mem_89_7_W0_clk),
    .W0_data(mem_89_7_W0_data),
    .W0_en(mem_89_7_W0_en),
    .W0_mask(mem_89_7_W0_mask)
  );
  split_mem_0_ext mem_90_0 (
    .R0_addr(mem_90_0_R0_addr),
    .R0_clk(mem_90_0_R0_clk),
    .R0_data(mem_90_0_R0_data),
    .R0_en(mem_90_0_R0_en),
    .W0_addr(mem_90_0_W0_addr),
    .W0_clk(mem_90_0_W0_clk),
    .W0_data(mem_90_0_W0_data),
    .W0_en(mem_90_0_W0_en),
    .W0_mask(mem_90_0_W0_mask)
  );
  split_mem_0_ext mem_90_1 (
    .R0_addr(mem_90_1_R0_addr),
    .R0_clk(mem_90_1_R0_clk),
    .R0_data(mem_90_1_R0_data),
    .R0_en(mem_90_1_R0_en),
    .W0_addr(mem_90_1_W0_addr),
    .W0_clk(mem_90_1_W0_clk),
    .W0_data(mem_90_1_W0_data),
    .W0_en(mem_90_1_W0_en),
    .W0_mask(mem_90_1_W0_mask)
  );
  split_mem_0_ext mem_90_2 (
    .R0_addr(mem_90_2_R0_addr),
    .R0_clk(mem_90_2_R0_clk),
    .R0_data(mem_90_2_R0_data),
    .R0_en(mem_90_2_R0_en),
    .W0_addr(mem_90_2_W0_addr),
    .W0_clk(mem_90_2_W0_clk),
    .W0_data(mem_90_2_W0_data),
    .W0_en(mem_90_2_W0_en),
    .W0_mask(mem_90_2_W0_mask)
  );
  split_mem_0_ext mem_90_3 (
    .R0_addr(mem_90_3_R0_addr),
    .R0_clk(mem_90_3_R0_clk),
    .R0_data(mem_90_3_R0_data),
    .R0_en(mem_90_3_R0_en),
    .W0_addr(mem_90_3_W0_addr),
    .W0_clk(mem_90_3_W0_clk),
    .W0_data(mem_90_3_W0_data),
    .W0_en(mem_90_3_W0_en),
    .W0_mask(mem_90_3_W0_mask)
  );
  split_mem_0_ext mem_90_4 (
    .R0_addr(mem_90_4_R0_addr),
    .R0_clk(mem_90_4_R0_clk),
    .R0_data(mem_90_4_R0_data),
    .R0_en(mem_90_4_R0_en),
    .W0_addr(mem_90_4_W0_addr),
    .W0_clk(mem_90_4_W0_clk),
    .W0_data(mem_90_4_W0_data),
    .W0_en(mem_90_4_W0_en),
    .W0_mask(mem_90_4_W0_mask)
  );
  split_mem_0_ext mem_90_5 (
    .R0_addr(mem_90_5_R0_addr),
    .R0_clk(mem_90_5_R0_clk),
    .R0_data(mem_90_5_R0_data),
    .R0_en(mem_90_5_R0_en),
    .W0_addr(mem_90_5_W0_addr),
    .W0_clk(mem_90_5_W0_clk),
    .W0_data(mem_90_5_W0_data),
    .W0_en(mem_90_5_W0_en),
    .W0_mask(mem_90_5_W0_mask)
  );
  split_mem_0_ext mem_90_6 (
    .R0_addr(mem_90_6_R0_addr),
    .R0_clk(mem_90_6_R0_clk),
    .R0_data(mem_90_6_R0_data),
    .R0_en(mem_90_6_R0_en),
    .W0_addr(mem_90_6_W0_addr),
    .W0_clk(mem_90_6_W0_clk),
    .W0_data(mem_90_6_W0_data),
    .W0_en(mem_90_6_W0_en),
    .W0_mask(mem_90_6_W0_mask)
  );
  split_mem_0_ext mem_90_7 (
    .R0_addr(mem_90_7_R0_addr),
    .R0_clk(mem_90_7_R0_clk),
    .R0_data(mem_90_7_R0_data),
    .R0_en(mem_90_7_R0_en),
    .W0_addr(mem_90_7_W0_addr),
    .W0_clk(mem_90_7_W0_clk),
    .W0_data(mem_90_7_W0_data),
    .W0_en(mem_90_7_W0_en),
    .W0_mask(mem_90_7_W0_mask)
  );
  split_mem_0_ext mem_91_0 (
    .R0_addr(mem_91_0_R0_addr),
    .R0_clk(mem_91_0_R0_clk),
    .R0_data(mem_91_0_R0_data),
    .R0_en(mem_91_0_R0_en),
    .W0_addr(mem_91_0_W0_addr),
    .W0_clk(mem_91_0_W0_clk),
    .W0_data(mem_91_0_W0_data),
    .W0_en(mem_91_0_W0_en),
    .W0_mask(mem_91_0_W0_mask)
  );
  split_mem_0_ext mem_91_1 (
    .R0_addr(mem_91_1_R0_addr),
    .R0_clk(mem_91_1_R0_clk),
    .R0_data(mem_91_1_R0_data),
    .R0_en(mem_91_1_R0_en),
    .W0_addr(mem_91_1_W0_addr),
    .W0_clk(mem_91_1_W0_clk),
    .W0_data(mem_91_1_W0_data),
    .W0_en(mem_91_1_W0_en),
    .W0_mask(mem_91_1_W0_mask)
  );
  split_mem_0_ext mem_91_2 (
    .R0_addr(mem_91_2_R0_addr),
    .R0_clk(mem_91_2_R0_clk),
    .R0_data(mem_91_2_R0_data),
    .R0_en(mem_91_2_R0_en),
    .W0_addr(mem_91_2_W0_addr),
    .W0_clk(mem_91_2_W0_clk),
    .W0_data(mem_91_2_W0_data),
    .W0_en(mem_91_2_W0_en),
    .W0_mask(mem_91_2_W0_mask)
  );
  split_mem_0_ext mem_91_3 (
    .R0_addr(mem_91_3_R0_addr),
    .R0_clk(mem_91_3_R0_clk),
    .R0_data(mem_91_3_R0_data),
    .R0_en(mem_91_3_R0_en),
    .W0_addr(mem_91_3_W0_addr),
    .W0_clk(mem_91_3_W0_clk),
    .W0_data(mem_91_3_W0_data),
    .W0_en(mem_91_3_W0_en),
    .W0_mask(mem_91_3_W0_mask)
  );
  split_mem_0_ext mem_91_4 (
    .R0_addr(mem_91_4_R0_addr),
    .R0_clk(mem_91_4_R0_clk),
    .R0_data(mem_91_4_R0_data),
    .R0_en(mem_91_4_R0_en),
    .W0_addr(mem_91_4_W0_addr),
    .W0_clk(mem_91_4_W0_clk),
    .W0_data(mem_91_4_W0_data),
    .W0_en(mem_91_4_W0_en),
    .W0_mask(mem_91_4_W0_mask)
  );
  split_mem_0_ext mem_91_5 (
    .R0_addr(mem_91_5_R0_addr),
    .R0_clk(mem_91_5_R0_clk),
    .R0_data(mem_91_5_R0_data),
    .R0_en(mem_91_5_R0_en),
    .W0_addr(mem_91_5_W0_addr),
    .W0_clk(mem_91_5_W0_clk),
    .W0_data(mem_91_5_W0_data),
    .W0_en(mem_91_5_W0_en),
    .W0_mask(mem_91_5_W0_mask)
  );
  split_mem_0_ext mem_91_6 (
    .R0_addr(mem_91_6_R0_addr),
    .R0_clk(mem_91_6_R0_clk),
    .R0_data(mem_91_6_R0_data),
    .R0_en(mem_91_6_R0_en),
    .W0_addr(mem_91_6_W0_addr),
    .W0_clk(mem_91_6_W0_clk),
    .W0_data(mem_91_6_W0_data),
    .W0_en(mem_91_6_W0_en),
    .W0_mask(mem_91_6_W0_mask)
  );
  split_mem_0_ext mem_91_7 (
    .R0_addr(mem_91_7_R0_addr),
    .R0_clk(mem_91_7_R0_clk),
    .R0_data(mem_91_7_R0_data),
    .R0_en(mem_91_7_R0_en),
    .W0_addr(mem_91_7_W0_addr),
    .W0_clk(mem_91_7_W0_clk),
    .W0_data(mem_91_7_W0_data),
    .W0_en(mem_91_7_W0_en),
    .W0_mask(mem_91_7_W0_mask)
  );
  split_mem_0_ext mem_92_0 (
    .R0_addr(mem_92_0_R0_addr),
    .R0_clk(mem_92_0_R0_clk),
    .R0_data(mem_92_0_R0_data),
    .R0_en(mem_92_0_R0_en),
    .W0_addr(mem_92_0_W0_addr),
    .W0_clk(mem_92_0_W0_clk),
    .W0_data(mem_92_0_W0_data),
    .W0_en(mem_92_0_W0_en),
    .W0_mask(mem_92_0_W0_mask)
  );
  split_mem_0_ext mem_92_1 (
    .R0_addr(mem_92_1_R0_addr),
    .R0_clk(mem_92_1_R0_clk),
    .R0_data(mem_92_1_R0_data),
    .R0_en(mem_92_1_R0_en),
    .W0_addr(mem_92_1_W0_addr),
    .W0_clk(mem_92_1_W0_clk),
    .W0_data(mem_92_1_W0_data),
    .W0_en(mem_92_1_W0_en),
    .W0_mask(mem_92_1_W0_mask)
  );
  split_mem_0_ext mem_92_2 (
    .R0_addr(mem_92_2_R0_addr),
    .R0_clk(mem_92_2_R0_clk),
    .R0_data(mem_92_2_R0_data),
    .R0_en(mem_92_2_R0_en),
    .W0_addr(mem_92_2_W0_addr),
    .W0_clk(mem_92_2_W0_clk),
    .W0_data(mem_92_2_W0_data),
    .W0_en(mem_92_2_W0_en),
    .W0_mask(mem_92_2_W0_mask)
  );
  split_mem_0_ext mem_92_3 (
    .R0_addr(mem_92_3_R0_addr),
    .R0_clk(mem_92_3_R0_clk),
    .R0_data(mem_92_3_R0_data),
    .R0_en(mem_92_3_R0_en),
    .W0_addr(mem_92_3_W0_addr),
    .W0_clk(mem_92_3_W0_clk),
    .W0_data(mem_92_3_W0_data),
    .W0_en(mem_92_3_W0_en),
    .W0_mask(mem_92_3_W0_mask)
  );
  split_mem_0_ext mem_92_4 (
    .R0_addr(mem_92_4_R0_addr),
    .R0_clk(mem_92_4_R0_clk),
    .R0_data(mem_92_4_R0_data),
    .R0_en(mem_92_4_R0_en),
    .W0_addr(mem_92_4_W0_addr),
    .W0_clk(mem_92_4_W0_clk),
    .W0_data(mem_92_4_W0_data),
    .W0_en(mem_92_4_W0_en),
    .W0_mask(mem_92_4_W0_mask)
  );
  split_mem_0_ext mem_92_5 (
    .R0_addr(mem_92_5_R0_addr),
    .R0_clk(mem_92_5_R0_clk),
    .R0_data(mem_92_5_R0_data),
    .R0_en(mem_92_5_R0_en),
    .W0_addr(mem_92_5_W0_addr),
    .W0_clk(mem_92_5_W0_clk),
    .W0_data(mem_92_5_W0_data),
    .W0_en(mem_92_5_W0_en),
    .W0_mask(mem_92_5_W0_mask)
  );
  split_mem_0_ext mem_92_6 (
    .R0_addr(mem_92_6_R0_addr),
    .R0_clk(mem_92_6_R0_clk),
    .R0_data(mem_92_6_R0_data),
    .R0_en(mem_92_6_R0_en),
    .W0_addr(mem_92_6_W0_addr),
    .W0_clk(mem_92_6_W0_clk),
    .W0_data(mem_92_6_W0_data),
    .W0_en(mem_92_6_W0_en),
    .W0_mask(mem_92_6_W0_mask)
  );
  split_mem_0_ext mem_92_7 (
    .R0_addr(mem_92_7_R0_addr),
    .R0_clk(mem_92_7_R0_clk),
    .R0_data(mem_92_7_R0_data),
    .R0_en(mem_92_7_R0_en),
    .W0_addr(mem_92_7_W0_addr),
    .W0_clk(mem_92_7_W0_clk),
    .W0_data(mem_92_7_W0_data),
    .W0_en(mem_92_7_W0_en),
    .W0_mask(mem_92_7_W0_mask)
  );
  split_mem_0_ext mem_93_0 (
    .R0_addr(mem_93_0_R0_addr),
    .R0_clk(mem_93_0_R0_clk),
    .R0_data(mem_93_0_R0_data),
    .R0_en(mem_93_0_R0_en),
    .W0_addr(mem_93_0_W0_addr),
    .W0_clk(mem_93_0_W0_clk),
    .W0_data(mem_93_0_W0_data),
    .W0_en(mem_93_0_W0_en),
    .W0_mask(mem_93_0_W0_mask)
  );
  split_mem_0_ext mem_93_1 (
    .R0_addr(mem_93_1_R0_addr),
    .R0_clk(mem_93_1_R0_clk),
    .R0_data(mem_93_1_R0_data),
    .R0_en(mem_93_1_R0_en),
    .W0_addr(mem_93_1_W0_addr),
    .W0_clk(mem_93_1_W0_clk),
    .W0_data(mem_93_1_W0_data),
    .W0_en(mem_93_1_W0_en),
    .W0_mask(mem_93_1_W0_mask)
  );
  split_mem_0_ext mem_93_2 (
    .R0_addr(mem_93_2_R0_addr),
    .R0_clk(mem_93_2_R0_clk),
    .R0_data(mem_93_2_R0_data),
    .R0_en(mem_93_2_R0_en),
    .W0_addr(mem_93_2_W0_addr),
    .W0_clk(mem_93_2_W0_clk),
    .W0_data(mem_93_2_W0_data),
    .W0_en(mem_93_2_W0_en),
    .W0_mask(mem_93_2_W0_mask)
  );
  split_mem_0_ext mem_93_3 (
    .R0_addr(mem_93_3_R0_addr),
    .R0_clk(mem_93_3_R0_clk),
    .R0_data(mem_93_3_R0_data),
    .R0_en(mem_93_3_R0_en),
    .W0_addr(mem_93_3_W0_addr),
    .W0_clk(mem_93_3_W0_clk),
    .W0_data(mem_93_3_W0_data),
    .W0_en(mem_93_3_W0_en),
    .W0_mask(mem_93_3_W0_mask)
  );
  split_mem_0_ext mem_93_4 (
    .R0_addr(mem_93_4_R0_addr),
    .R0_clk(mem_93_4_R0_clk),
    .R0_data(mem_93_4_R0_data),
    .R0_en(mem_93_4_R0_en),
    .W0_addr(mem_93_4_W0_addr),
    .W0_clk(mem_93_4_W0_clk),
    .W0_data(mem_93_4_W0_data),
    .W0_en(mem_93_4_W0_en),
    .W0_mask(mem_93_4_W0_mask)
  );
  split_mem_0_ext mem_93_5 (
    .R0_addr(mem_93_5_R0_addr),
    .R0_clk(mem_93_5_R0_clk),
    .R0_data(mem_93_5_R0_data),
    .R0_en(mem_93_5_R0_en),
    .W0_addr(mem_93_5_W0_addr),
    .W0_clk(mem_93_5_W0_clk),
    .W0_data(mem_93_5_W0_data),
    .W0_en(mem_93_5_W0_en),
    .W0_mask(mem_93_5_W0_mask)
  );
  split_mem_0_ext mem_93_6 (
    .R0_addr(mem_93_6_R0_addr),
    .R0_clk(mem_93_6_R0_clk),
    .R0_data(mem_93_6_R0_data),
    .R0_en(mem_93_6_R0_en),
    .W0_addr(mem_93_6_W0_addr),
    .W0_clk(mem_93_6_W0_clk),
    .W0_data(mem_93_6_W0_data),
    .W0_en(mem_93_6_W0_en),
    .W0_mask(mem_93_6_W0_mask)
  );
  split_mem_0_ext mem_93_7 (
    .R0_addr(mem_93_7_R0_addr),
    .R0_clk(mem_93_7_R0_clk),
    .R0_data(mem_93_7_R0_data),
    .R0_en(mem_93_7_R0_en),
    .W0_addr(mem_93_7_W0_addr),
    .W0_clk(mem_93_7_W0_clk),
    .W0_data(mem_93_7_W0_data),
    .W0_en(mem_93_7_W0_en),
    .W0_mask(mem_93_7_W0_mask)
  );
  split_mem_0_ext mem_94_0 (
    .R0_addr(mem_94_0_R0_addr),
    .R0_clk(mem_94_0_R0_clk),
    .R0_data(mem_94_0_R0_data),
    .R0_en(mem_94_0_R0_en),
    .W0_addr(mem_94_0_W0_addr),
    .W0_clk(mem_94_0_W0_clk),
    .W0_data(mem_94_0_W0_data),
    .W0_en(mem_94_0_W0_en),
    .W0_mask(mem_94_0_W0_mask)
  );
  split_mem_0_ext mem_94_1 (
    .R0_addr(mem_94_1_R0_addr),
    .R0_clk(mem_94_1_R0_clk),
    .R0_data(mem_94_1_R0_data),
    .R0_en(mem_94_1_R0_en),
    .W0_addr(mem_94_1_W0_addr),
    .W0_clk(mem_94_1_W0_clk),
    .W0_data(mem_94_1_W0_data),
    .W0_en(mem_94_1_W0_en),
    .W0_mask(mem_94_1_W0_mask)
  );
  split_mem_0_ext mem_94_2 (
    .R0_addr(mem_94_2_R0_addr),
    .R0_clk(mem_94_2_R0_clk),
    .R0_data(mem_94_2_R0_data),
    .R0_en(mem_94_2_R0_en),
    .W0_addr(mem_94_2_W0_addr),
    .W0_clk(mem_94_2_W0_clk),
    .W0_data(mem_94_2_W0_data),
    .W0_en(mem_94_2_W0_en),
    .W0_mask(mem_94_2_W0_mask)
  );
  split_mem_0_ext mem_94_3 (
    .R0_addr(mem_94_3_R0_addr),
    .R0_clk(mem_94_3_R0_clk),
    .R0_data(mem_94_3_R0_data),
    .R0_en(mem_94_3_R0_en),
    .W0_addr(mem_94_3_W0_addr),
    .W0_clk(mem_94_3_W0_clk),
    .W0_data(mem_94_3_W0_data),
    .W0_en(mem_94_3_W0_en),
    .W0_mask(mem_94_3_W0_mask)
  );
  split_mem_0_ext mem_94_4 (
    .R0_addr(mem_94_4_R0_addr),
    .R0_clk(mem_94_4_R0_clk),
    .R0_data(mem_94_4_R0_data),
    .R0_en(mem_94_4_R0_en),
    .W0_addr(mem_94_4_W0_addr),
    .W0_clk(mem_94_4_W0_clk),
    .W0_data(mem_94_4_W0_data),
    .W0_en(mem_94_4_W0_en),
    .W0_mask(mem_94_4_W0_mask)
  );
  split_mem_0_ext mem_94_5 (
    .R0_addr(mem_94_5_R0_addr),
    .R0_clk(mem_94_5_R0_clk),
    .R0_data(mem_94_5_R0_data),
    .R0_en(mem_94_5_R0_en),
    .W0_addr(mem_94_5_W0_addr),
    .W0_clk(mem_94_5_W0_clk),
    .W0_data(mem_94_5_W0_data),
    .W0_en(mem_94_5_W0_en),
    .W0_mask(mem_94_5_W0_mask)
  );
  split_mem_0_ext mem_94_6 (
    .R0_addr(mem_94_6_R0_addr),
    .R0_clk(mem_94_6_R0_clk),
    .R0_data(mem_94_6_R0_data),
    .R0_en(mem_94_6_R0_en),
    .W0_addr(mem_94_6_W0_addr),
    .W0_clk(mem_94_6_W0_clk),
    .W0_data(mem_94_6_W0_data),
    .W0_en(mem_94_6_W0_en),
    .W0_mask(mem_94_6_W0_mask)
  );
  split_mem_0_ext mem_94_7 (
    .R0_addr(mem_94_7_R0_addr),
    .R0_clk(mem_94_7_R0_clk),
    .R0_data(mem_94_7_R0_data),
    .R0_en(mem_94_7_R0_en),
    .W0_addr(mem_94_7_W0_addr),
    .W0_clk(mem_94_7_W0_clk),
    .W0_data(mem_94_7_W0_data),
    .W0_en(mem_94_7_W0_en),
    .W0_mask(mem_94_7_W0_mask)
  );
  split_mem_0_ext mem_95_0 (
    .R0_addr(mem_95_0_R0_addr),
    .R0_clk(mem_95_0_R0_clk),
    .R0_data(mem_95_0_R0_data),
    .R0_en(mem_95_0_R0_en),
    .W0_addr(mem_95_0_W0_addr),
    .W0_clk(mem_95_0_W0_clk),
    .W0_data(mem_95_0_W0_data),
    .W0_en(mem_95_0_W0_en),
    .W0_mask(mem_95_0_W0_mask)
  );
  split_mem_0_ext mem_95_1 (
    .R0_addr(mem_95_1_R0_addr),
    .R0_clk(mem_95_1_R0_clk),
    .R0_data(mem_95_1_R0_data),
    .R0_en(mem_95_1_R0_en),
    .W0_addr(mem_95_1_W0_addr),
    .W0_clk(mem_95_1_W0_clk),
    .W0_data(mem_95_1_W0_data),
    .W0_en(mem_95_1_W0_en),
    .W0_mask(mem_95_1_W0_mask)
  );
  split_mem_0_ext mem_95_2 (
    .R0_addr(mem_95_2_R0_addr),
    .R0_clk(mem_95_2_R0_clk),
    .R0_data(mem_95_2_R0_data),
    .R0_en(mem_95_2_R0_en),
    .W0_addr(mem_95_2_W0_addr),
    .W0_clk(mem_95_2_W0_clk),
    .W0_data(mem_95_2_W0_data),
    .W0_en(mem_95_2_W0_en),
    .W0_mask(mem_95_2_W0_mask)
  );
  split_mem_0_ext mem_95_3 (
    .R0_addr(mem_95_3_R0_addr),
    .R0_clk(mem_95_3_R0_clk),
    .R0_data(mem_95_3_R0_data),
    .R0_en(mem_95_3_R0_en),
    .W0_addr(mem_95_3_W0_addr),
    .W0_clk(mem_95_3_W0_clk),
    .W0_data(mem_95_3_W0_data),
    .W0_en(mem_95_3_W0_en),
    .W0_mask(mem_95_3_W0_mask)
  );
  split_mem_0_ext mem_95_4 (
    .R0_addr(mem_95_4_R0_addr),
    .R0_clk(mem_95_4_R0_clk),
    .R0_data(mem_95_4_R0_data),
    .R0_en(mem_95_4_R0_en),
    .W0_addr(mem_95_4_W0_addr),
    .W0_clk(mem_95_4_W0_clk),
    .W0_data(mem_95_4_W0_data),
    .W0_en(mem_95_4_W0_en),
    .W0_mask(mem_95_4_W0_mask)
  );
  split_mem_0_ext mem_95_5 (
    .R0_addr(mem_95_5_R0_addr),
    .R0_clk(mem_95_5_R0_clk),
    .R0_data(mem_95_5_R0_data),
    .R0_en(mem_95_5_R0_en),
    .W0_addr(mem_95_5_W0_addr),
    .W0_clk(mem_95_5_W0_clk),
    .W0_data(mem_95_5_W0_data),
    .W0_en(mem_95_5_W0_en),
    .W0_mask(mem_95_5_W0_mask)
  );
  split_mem_0_ext mem_95_6 (
    .R0_addr(mem_95_6_R0_addr),
    .R0_clk(mem_95_6_R0_clk),
    .R0_data(mem_95_6_R0_data),
    .R0_en(mem_95_6_R0_en),
    .W0_addr(mem_95_6_W0_addr),
    .W0_clk(mem_95_6_W0_clk),
    .W0_data(mem_95_6_W0_data),
    .W0_en(mem_95_6_W0_en),
    .W0_mask(mem_95_6_W0_mask)
  );
  split_mem_0_ext mem_95_7 (
    .R0_addr(mem_95_7_R0_addr),
    .R0_clk(mem_95_7_R0_clk),
    .R0_data(mem_95_7_R0_data),
    .R0_en(mem_95_7_R0_en),
    .W0_addr(mem_95_7_W0_addr),
    .W0_clk(mem_95_7_W0_clk),
    .W0_data(mem_95_7_W0_data),
    .W0_en(mem_95_7_W0_en),
    .W0_mask(mem_95_7_W0_mask)
  );
  split_mem_0_ext mem_96_0 (
    .R0_addr(mem_96_0_R0_addr),
    .R0_clk(mem_96_0_R0_clk),
    .R0_data(mem_96_0_R0_data),
    .R0_en(mem_96_0_R0_en),
    .W0_addr(mem_96_0_W0_addr),
    .W0_clk(mem_96_0_W0_clk),
    .W0_data(mem_96_0_W0_data),
    .W0_en(mem_96_0_W0_en),
    .W0_mask(mem_96_0_W0_mask)
  );
  split_mem_0_ext mem_96_1 (
    .R0_addr(mem_96_1_R0_addr),
    .R0_clk(mem_96_1_R0_clk),
    .R0_data(mem_96_1_R0_data),
    .R0_en(mem_96_1_R0_en),
    .W0_addr(mem_96_1_W0_addr),
    .W0_clk(mem_96_1_W0_clk),
    .W0_data(mem_96_1_W0_data),
    .W0_en(mem_96_1_W0_en),
    .W0_mask(mem_96_1_W0_mask)
  );
  split_mem_0_ext mem_96_2 (
    .R0_addr(mem_96_2_R0_addr),
    .R0_clk(mem_96_2_R0_clk),
    .R0_data(mem_96_2_R0_data),
    .R0_en(mem_96_2_R0_en),
    .W0_addr(mem_96_2_W0_addr),
    .W0_clk(mem_96_2_W0_clk),
    .W0_data(mem_96_2_W0_data),
    .W0_en(mem_96_2_W0_en),
    .W0_mask(mem_96_2_W0_mask)
  );
  split_mem_0_ext mem_96_3 (
    .R0_addr(mem_96_3_R0_addr),
    .R0_clk(mem_96_3_R0_clk),
    .R0_data(mem_96_3_R0_data),
    .R0_en(mem_96_3_R0_en),
    .W0_addr(mem_96_3_W0_addr),
    .W0_clk(mem_96_3_W0_clk),
    .W0_data(mem_96_3_W0_data),
    .W0_en(mem_96_3_W0_en),
    .W0_mask(mem_96_3_W0_mask)
  );
  split_mem_0_ext mem_96_4 (
    .R0_addr(mem_96_4_R0_addr),
    .R0_clk(mem_96_4_R0_clk),
    .R0_data(mem_96_4_R0_data),
    .R0_en(mem_96_4_R0_en),
    .W0_addr(mem_96_4_W0_addr),
    .W0_clk(mem_96_4_W0_clk),
    .W0_data(mem_96_4_W0_data),
    .W0_en(mem_96_4_W0_en),
    .W0_mask(mem_96_4_W0_mask)
  );
  split_mem_0_ext mem_96_5 (
    .R0_addr(mem_96_5_R0_addr),
    .R0_clk(mem_96_5_R0_clk),
    .R0_data(mem_96_5_R0_data),
    .R0_en(mem_96_5_R0_en),
    .W0_addr(mem_96_5_W0_addr),
    .W0_clk(mem_96_5_W0_clk),
    .W0_data(mem_96_5_W0_data),
    .W0_en(mem_96_5_W0_en),
    .W0_mask(mem_96_5_W0_mask)
  );
  split_mem_0_ext mem_96_6 (
    .R0_addr(mem_96_6_R0_addr),
    .R0_clk(mem_96_6_R0_clk),
    .R0_data(mem_96_6_R0_data),
    .R0_en(mem_96_6_R0_en),
    .W0_addr(mem_96_6_W0_addr),
    .W0_clk(mem_96_6_W0_clk),
    .W0_data(mem_96_6_W0_data),
    .W0_en(mem_96_6_W0_en),
    .W0_mask(mem_96_6_W0_mask)
  );
  split_mem_0_ext mem_96_7 (
    .R0_addr(mem_96_7_R0_addr),
    .R0_clk(mem_96_7_R0_clk),
    .R0_data(mem_96_7_R0_data),
    .R0_en(mem_96_7_R0_en),
    .W0_addr(mem_96_7_W0_addr),
    .W0_clk(mem_96_7_W0_clk),
    .W0_data(mem_96_7_W0_data),
    .W0_en(mem_96_7_W0_en),
    .W0_mask(mem_96_7_W0_mask)
  );
  split_mem_0_ext mem_97_0 (
    .R0_addr(mem_97_0_R0_addr),
    .R0_clk(mem_97_0_R0_clk),
    .R0_data(mem_97_0_R0_data),
    .R0_en(mem_97_0_R0_en),
    .W0_addr(mem_97_0_W0_addr),
    .W0_clk(mem_97_0_W0_clk),
    .W0_data(mem_97_0_W0_data),
    .W0_en(mem_97_0_W0_en),
    .W0_mask(mem_97_0_W0_mask)
  );
  split_mem_0_ext mem_97_1 (
    .R0_addr(mem_97_1_R0_addr),
    .R0_clk(mem_97_1_R0_clk),
    .R0_data(mem_97_1_R0_data),
    .R0_en(mem_97_1_R0_en),
    .W0_addr(mem_97_1_W0_addr),
    .W0_clk(mem_97_1_W0_clk),
    .W0_data(mem_97_1_W0_data),
    .W0_en(mem_97_1_W0_en),
    .W0_mask(mem_97_1_W0_mask)
  );
  split_mem_0_ext mem_97_2 (
    .R0_addr(mem_97_2_R0_addr),
    .R0_clk(mem_97_2_R0_clk),
    .R0_data(mem_97_2_R0_data),
    .R0_en(mem_97_2_R0_en),
    .W0_addr(mem_97_2_W0_addr),
    .W0_clk(mem_97_2_W0_clk),
    .W0_data(mem_97_2_W0_data),
    .W0_en(mem_97_2_W0_en),
    .W0_mask(mem_97_2_W0_mask)
  );
  split_mem_0_ext mem_97_3 (
    .R0_addr(mem_97_3_R0_addr),
    .R0_clk(mem_97_3_R0_clk),
    .R0_data(mem_97_3_R0_data),
    .R0_en(mem_97_3_R0_en),
    .W0_addr(mem_97_3_W0_addr),
    .W0_clk(mem_97_3_W0_clk),
    .W0_data(mem_97_3_W0_data),
    .W0_en(mem_97_3_W0_en),
    .W0_mask(mem_97_3_W0_mask)
  );
  split_mem_0_ext mem_97_4 (
    .R0_addr(mem_97_4_R0_addr),
    .R0_clk(mem_97_4_R0_clk),
    .R0_data(mem_97_4_R0_data),
    .R0_en(mem_97_4_R0_en),
    .W0_addr(mem_97_4_W0_addr),
    .W0_clk(mem_97_4_W0_clk),
    .W0_data(mem_97_4_W0_data),
    .W0_en(mem_97_4_W0_en),
    .W0_mask(mem_97_4_W0_mask)
  );
  split_mem_0_ext mem_97_5 (
    .R0_addr(mem_97_5_R0_addr),
    .R0_clk(mem_97_5_R0_clk),
    .R0_data(mem_97_5_R0_data),
    .R0_en(mem_97_5_R0_en),
    .W0_addr(mem_97_5_W0_addr),
    .W0_clk(mem_97_5_W0_clk),
    .W0_data(mem_97_5_W0_data),
    .W0_en(mem_97_5_W0_en),
    .W0_mask(mem_97_5_W0_mask)
  );
  split_mem_0_ext mem_97_6 (
    .R0_addr(mem_97_6_R0_addr),
    .R0_clk(mem_97_6_R0_clk),
    .R0_data(mem_97_6_R0_data),
    .R0_en(mem_97_6_R0_en),
    .W0_addr(mem_97_6_W0_addr),
    .W0_clk(mem_97_6_W0_clk),
    .W0_data(mem_97_6_W0_data),
    .W0_en(mem_97_6_W0_en),
    .W0_mask(mem_97_6_W0_mask)
  );
  split_mem_0_ext mem_97_7 (
    .R0_addr(mem_97_7_R0_addr),
    .R0_clk(mem_97_7_R0_clk),
    .R0_data(mem_97_7_R0_data),
    .R0_en(mem_97_7_R0_en),
    .W0_addr(mem_97_7_W0_addr),
    .W0_clk(mem_97_7_W0_clk),
    .W0_data(mem_97_7_W0_data),
    .W0_en(mem_97_7_W0_en),
    .W0_mask(mem_97_7_W0_mask)
  );
  split_mem_0_ext mem_98_0 (
    .R0_addr(mem_98_0_R0_addr),
    .R0_clk(mem_98_0_R0_clk),
    .R0_data(mem_98_0_R0_data),
    .R0_en(mem_98_0_R0_en),
    .W0_addr(mem_98_0_W0_addr),
    .W0_clk(mem_98_0_W0_clk),
    .W0_data(mem_98_0_W0_data),
    .W0_en(mem_98_0_W0_en),
    .W0_mask(mem_98_0_W0_mask)
  );
  split_mem_0_ext mem_98_1 (
    .R0_addr(mem_98_1_R0_addr),
    .R0_clk(mem_98_1_R0_clk),
    .R0_data(mem_98_1_R0_data),
    .R0_en(mem_98_1_R0_en),
    .W0_addr(mem_98_1_W0_addr),
    .W0_clk(mem_98_1_W0_clk),
    .W0_data(mem_98_1_W0_data),
    .W0_en(mem_98_1_W0_en),
    .W0_mask(mem_98_1_W0_mask)
  );
  split_mem_0_ext mem_98_2 (
    .R0_addr(mem_98_2_R0_addr),
    .R0_clk(mem_98_2_R0_clk),
    .R0_data(mem_98_2_R0_data),
    .R0_en(mem_98_2_R0_en),
    .W0_addr(mem_98_2_W0_addr),
    .W0_clk(mem_98_2_W0_clk),
    .W0_data(mem_98_2_W0_data),
    .W0_en(mem_98_2_W0_en),
    .W0_mask(mem_98_2_W0_mask)
  );
  split_mem_0_ext mem_98_3 (
    .R0_addr(mem_98_3_R0_addr),
    .R0_clk(mem_98_3_R0_clk),
    .R0_data(mem_98_3_R0_data),
    .R0_en(mem_98_3_R0_en),
    .W0_addr(mem_98_3_W0_addr),
    .W0_clk(mem_98_3_W0_clk),
    .W0_data(mem_98_3_W0_data),
    .W0_en(mem_98_3_W0_en),
    .W0_mask(mem_98_3_W0_mask)
  );
  split_mem_0_ext mem_98_4 (
    .R0_addr(mem_98_4_R0_addr),
    .R0_clk(mem_98_4_R0_clk),
    .R0_data(mem_98_4_R0_data),
    .R0_en(mem_98_4_R0_en),
    .W0_addr(mem_98_4_W0_addr),
    .W0_clk(mem_98_4_W0_clk),
    .W0_data(mem_98_4_W0_data),
    .W0_en(mem_98_4_W0_en),
    .W0_mask(mem_98_4_W0_mask)
  );
  split_mem_0_ext mem_98_5 (
    .R0_addr(mem_98_5_R0_addr),
    .R0_clk(mem_98_5_R0_clk),
    .R0_data(mem_98_5_R0_data),
    .R0_en(mem_98_5_R0_en),
    .W0_addr(mem_98_5_W0_addr),
    .W0_clk(mem_98_5_W0_clk),
    .W0_data(mem_98_5_W0_data),
    .W0_en(mem_98_5_W0_en),
    .W0_mask(mem_98_5_W0_mask)
  );
  split_mem_0_ext mem_98_6 (
    .R0_addr(mem_98_6_R0_addr),
    .R0_clk(mem_98_6_R0_clk),
    .R0_data(mem_98_6_R0_data),
    .R0_en(mem_98_6_R0_en),
    .W0_addr(mem_98_6_W0_addr),
    .W0_clk(mem_98_6_W0_clk),
    .W0_data(mem_98_6_W0_data),
    .W0_en(mem_98_6_W0_en),
    .W0_mask(mem_98_6_W0_mask)
  );
  split_mem_0_ext mem_98_7 (
    .R0_addr(mem_98_7_R0_addr),
    .R0_clk(mem_98_7_R0_clk),
    .R0_data(mem_98_7_R0_data),
    .R0_en(mem_98_7_R0_en),
    .W0_addr(mem_98_7_W0_addr),
    .W0_clk(mem_98_7_W0_clk),
    .W0_data(mem_98_7_W0_data),
    .W0_en(mem_98_7_W0_en),
    .W0_mask(mem_98_7_W0_mask)
  );
  split_mem_0_ext mem_99_0 (
    .R0_addr(mem_99_0_R0_addr),
    .R0_clk(mem_99_0_R0_clk),
    .R0_data(mem_99_0_R0_data),
    .R0_en(mem_99_0_R0_en),
    .W0_addr(mem_99_0_W0_addr),
    .W0_clk(mem_99_0_W0_clk),
    .W0_data(mem_99_0_W0_data),
    .W0_en(mem_99_0_W0_en),
    .W0_mask(mem_99_0_W0_mask)
  );
  split_mem_0_ext mem_99_1 (
    .R0_addr(mem_99_1_R0_addr),
    .R0_clk(mem_99_1_R0_clk),
    .R0_data(mem_99_1_R0_data),
    .R0_en(mem_99_1_R0_en),
    .W0_addr(mem_99_1_W0_addr),
    .W0_clk(mem_99_1_W0_clk),
    .W0_data(mem_99_1_W0_data),
    .W0_en(mem_99_1_W0_en),
    .W0_mask(mem_99_1_W0_mask)
  );
  split_mem_0_ext mem_99_2 (
    .R0_addr(mem_99_2_R0_addr),
    .R0_clk(mem_99_2_R0_clk),
    .R0_data(mem_99_2_R0_data),
    .R0_en(mem_99_2_R0_en),
    .W0_addr(mem_99_2_W0_addr),
    .W0_clk(mem_99_2_W0_clk),
    .W0_data(mem_99_2_W0_data),
    .W0_en(mem_99_2_W0_en),
    .W0_mask(mem_99_2_W0_mask)
  );
  split_mem_0_ext mem_99_3 (
    .R0_addr(mem_99_3_R0_addr),
    .R0_clk(mem_99_3_R0_clk),
    .R0_data(mem_99_3_R0_data),
    .R0_en(mem_99_3_R0_en),
    .W0_addr(mem_99_3_W0_addr),
    .W0_clk(mem_99_3_W0_clk),
    .W0_data(mem_99_3_W0_data),
    .W0_en(mem_99_3_W0_en),
    .W0_mask(mem_99_3_W0_mask)
  );
  split_mem_0_ext mem_99_4 (
    .R0_addr(mem_99_4_R0_addr),
    .R0_clk(mem_99_4_R0_clk),
    .R0_data(mem_99_4_R0_data),
    .R0_en(mem_99_4_R0_en),
    .W0_addr(mem_99_4_W0_addr),
    .W0_clk(mem_99_4_W0_clk),
    .W0_data(mem_99_4_W0_data),
    .W0_en(mem_99_4_W0_en),
    .W0_mask(mem_99_4_W0_mask)
  );
  split_mem_0_ext mem_99_5 (
    .R0_addr(mem_99_5_R0_addr),
    .R0_clk(mem_99_5_R0_clk),
    .R0_data(mem_99_5_R0_data),
    .R0_en(mem_99_5_R0_en),
    .W0_addr(mem_99_5_W0_addr),
    .W0_clk(mem_99_5_W0_clk),
    .W0_data(mem_99_5_W0_data),
    .W0_en(mem_99_5_W0_en),
    .W0_mask(mem_99_5_W0_mask)
  );
  split_mem_0_ext mem_99_6 (
    .R0_addr(mem_99_6_R0_addr),
    .R0_clk(mem_99_6_R0_clk),
    .R0_data(mem_99_6_R0_data),
    .R0_en(mem_99_6_R0_en),
    .W0_addr(mem_99_6_W0_addr),
    .W0_clk(mem_99_6_W0_clk),
    .W0_data(mem_99_6_W0_data),
    .W0_en(mem_99_6_W0_en),
    .W0_mask(mem_99_6_W0_mask)
  );
  split_mem_0_ext mem_99_7 (
    .R0_addr(mem_99_7_R0_addr),
    .R0_clk(mem_99_7_R0_clk),
    .R0_data(mem_99_7_R0_data),
    .R0_en(mem_99_7_R0_en),
    .W0_addr(mem_99_7_W0_addr),
    .W0_clk(mem_99_7_W0_clk),
    .W0_data(mem_99_7_W0_data),
    .W0_en(mem_99_7_W0_en),
    .W0_mask(mem_99_7_W0_mask)
  );
  split_mem_0_ext mem_100_0 (
    .R0_addr(mem_100_0_R0_addr),
    .R0_clk(mem_100_0_R0_clk),
    .R0_data(mem_100_0_R0_data),
    .R0_en(mem_100_0_R0_en),
    .W0_addr(mem_100_0_W0_addr),
    .W0_clk(mem_100_0_W0_clk),
    .W0_data(mem_100_0_W0_data),
    .W0_en(mem_100_0_W0_en),
    .W0_mask(mem_100_0_W0_mask)
  );
  split_mem_0_ext mem_100_1 (
    .R0_addr(mem_100_1_R0_addr),
    .R0_clk(mem_100_1_R0_clk),
    .R0_data(mem_100_1_R0_data),
    .R0_en(mem_100_1_R0_en),
    .W0_addr(mem_100_1_W0_addr),
    .W0_clk(mem_100_1_W0_clk),
    .W0_data(mem_100_1_W0_data),
    .W0_en(mem_100_1_W0_en),
    .W0_mask(mem_100_1_W0_mask)
  );
  split_mem_0_ext mem_100_2 (
    .R0_addr(mem_100_2_R0_addr),
    .R0_clk(mem_100_2_R0_clk),
    .R0_data(mem_100_2_R0_data),
    .R0_en(mem_100_2_R0_en),
    .W0_addr(mem_100_2_W0_addr),
    .W0_clk(mem_100_2_W0_clk),
    .W0_data(mem_100_2_W0_data),
    .W0_en(mem_100_2_W0_en),
    .W0_mask(mem_100_2_W0_mask)
  );
  split_mem_0_ext mem_100_3 (
    .R0_addr(mem_100_3_R0_addr),
    .R0_clk(mem_100_3_R0_clk),
    .R0_data(mem_100_3_R0_data),
    .R0_en(mem_100_3_R0_en),
    .W0_addr(mem_100_3_W0_addr),
    .W0_clk(mem_100_3_W0_clk),
    .W0_data(mem_100_3_W0_data),
    .W0_en(mem_100_3_W0_en),
    .W0_mask(mem_100_3_W0_mask)
  );
  split_mem_0_ext mem_100_4 (
    .R0_addr(mem_100_4_R0_addr),
    .R0_clk(mem_100_4_R0_clk),
    .R0_data(mem_100_4_R0_data),
    .R0_en(mem_100_4_R0_en),
    .W0_addr(mem_100_4_W0_addr),
    .W0_clk(mem_100_4_W0_clk),
    .W0_data(mem_100_4_W0_data),
    .W0_en(mem_100_4_W0_en),
    .W0_mask(mem_100_4_W0_mask)
  );
  split_mem_0_ext mem_100_5 (
    .R0_addr(mem_100_5_R0_addr),
    .R0_clk(mem_100_5_R0_clk),
    .R0_data(mem_100_5_R0_data),
    .R0_en(mem_100_5_R0_en),
    .W0_addr(mem_100_5_W0_addr),
    .W0_clk(mem_100_5_W0_clk),
    .W0_data(mem_100_5_W0_data),
    .W0_en(mem_100_5_W0_en),
    .W0_mask(mem_100_5_W0_mask)
  );
  split_mem_0_ext mem_100_6 (
    .R0_addr(mem_100_6_R0_addr),
    .R0_clk(mem_100_6_R0_clk),
    .R0_data(mem_100_6_R0_data),
    .R0_en(mem_100_6_R0_en),
    .W0_addr(mem_100_6_W0_addr),
    .W0_clk(mem_100_6_W0_clk),
    .W0_data(mem_100_6_W0_data),
    .W0_en(mem_100_6_W0_en),
    .W0_mask(mem_100_6_W0_mask)
  );
  split_mem_0_ext mem_100_7 (
    .R0_addr(mem_100_7_R0_addr),
    .R0_clk(mem_100_7_R0_clk),
    .R0_data(mem_100_7_R0_data),
    .R0_en(mem_100_7_R0_en),
    .W0_addr(mem_100_7_W0_addr),
    .W0_clk(mem_100_7_W0_clk),
    .W0_data(mem_100_7_W0_data),
    .W0_en(mem_100_7_W0_en),
    .W0_mask(mem_100_7_W0_mask)
  );
  split_mem_0_ext mem_101_0 (
    .R0_addr(mem_101_0_R0_addr),
    .R0_clk(mem_101_0_R0_clk),
    .R0_data(mem_101_0_R0_data),
    .R0_en(mem_101_0_R0_en),
    .W0_addr(mem_101_0_W0_addr),
    .W0_clk(mem_101_0_W0_clk),
    .W0_data(mem_101_0_W0_data),
    .W0_en(mem_101_0_W0_en),
    .W0_mask(mem_101_0_W0_mask)
  );
  split_mem_0_ext mem_101_1 (
    .R0_addr(mem_101_1_R0_addr),
    .R0_clk(mem_101_1_R0_clk),
    .R0_data(mem_101_1_R0_data),
    .R0_en(mem_101_1_R0_en),
    .W0_addr(mem_101_1_W0_addr),
    .W0_clk(mem_101_1_W0_clk),
    .W0_data(mem_101_1_W0_data),
    .W0_en(mem_101_1_W0_en),
    .W0_mask(mem_101_1_W0_mask)
  );
  split_mem_0_ext mem_101_2 (
    .R0_addr(mem_101_2_R0_addr),
    .R0_clk(mem_101_2_R0_clk),
    .R0_data(mem_101_2_R0_data),
    .R0_en(mem_101_2_R0_en),
    .W0_addr(mem_101_2_W0_addr),
    .W0_clk(mem_101_2_W0_clk),
    .W0_data(mem_101_2_W0_data),
    .W0_en(mem_101_2_W0_en),
    .W0_mask(mem_101_2_W0_mask)
  );
  split_mem_0_ext mem_101_3 (
    .R0_addr(mem_101_3_R0_addr),
    .R0_clk(mem_101_3_R0_clk),
    .R0_data(mem_101_3_R0_data),
    .R0_en(mem_101_3_R0_en),
    .W0_addr(mem_101_3_W0_addr),
    .W0_clk(mem_101_3_W0_clk),
    .W0_data(mem_101_3_W0_data),
    .W0_en(mem_101_3_W0_en),
    .W0_mask(mem_101_3_W0_mask)
  );
  split_mem_0_ext mem_101_4 (
    .R0_addr(mem_101_4_R0_addr),
    .R0_clk(mem_101_4_R0_clk),
    .R0_data(mem_101_4_R0_data),
    .R0_en(mem_101_4_R0_en),
    .W0_addr(mem_101_4_W0_addr),
    .W0_clk(mem_101_4_W0_clk),
    .W0_data(mem_101_4_W0_data),
    .W0_en(mem_101_4_W0_en),
    .W0_mask(mem_101_4_W0_mask)
  );
  split_mem_0_ext mem_101_5 (
    .R0_addr(mem_101_5_R0_addr),
    .R0_clk(mem_101_5_R0_clk),
    .R0_data(mem_101_5_R0_data),
    .R0_en(mem_101_5_R0_en),
    .W0_addr(mem_101_5_W0_addr),
    .W0_clk(mem_101_5_W0_clk),
    .W0_data(mem_101_5_W0_data),
    .W0_en(mem_101_5_W0_en),
    .W0_mask(mem_101_5_W0_mask)
  );
  split_mem_0_ext mem_101_6 (
    .R0_addr(mem_101_6_R0_addr),
    .R0_clk(mem_101_6_R0_clk),
    .R0_data(mem_101_6_R0_data),
    .R0_en(mem_101_6_R0_en),
    .W0_addr(mem_101_6_W0_addr),
    .W0_clk(mem_101_6_W0_clk),
    .W0_data(mem_101_6_W0_data),
    .W0_en(mem_101_6_W0_en),
    .W0_mask(mem_101_6_W0_mask)
  );
  split_mem_0_ext mem_101_7 (
    .R0_addr(mem_101_7_R0_addr),
    .R0_clk(mem_101_7_R0_clk),
    .R0_data(mem_101_7_R0_data),
    .R0_en(mem_101_7_R0_en),
    .W0_addr(mem_101_7_W0_addr),
    .W0_clk(mem_101_7_W0_clk),
    .W0_data(mem_101_7_W0_data),
    .W0_en(mem_101_7_W0_en),
    .W0_mask(mem_101_7_W0_mask)
  );
  split_mem_0_ext mem_102_0 (
    .R0_addr(mem_102_0_R0_addr),
    .R0_clk(mem_102_0_R0_clk),
    .R0_data(mem_102_0_R0_data),
    .R0_en(mem_102_0_R0_en),
    .W0_addr(mem_102_0_W0_addr),
    .W0_clk(mem_102_0_W0_clk),
    .W0_data(mem_102_0_W0_data),
    .W0_en(mem_102_0_W0_en),
    .W0_mask(mem_102_0_W0_mask)
  );
  split_mem_0_ext mem_102_1 (
    .R0_addr(mem_102_1_R0_addr),
    .R0_clk(mem_102_1_R0_clk),
    .R0_data(mem_102_1_R0_data),
    .R0_en(mem_102_1_R0_en),
    .W0_addr(mem_102_1_W0_addr),
    .W0_clk(mem_102_1_W0_clk),
    .W0_data(mem_102_1_W0_data),
    .W0_en(mem_102_1_W0_en),
    .W0_mask(mem_102_1_W0_mask)
  );
  split_mem_0_ext mem_102_2 (
    .R0_addr(mem_102_2_R0_addr),
    .R0_clk(mem_102_2_R0_clk),
    .R0_data(mem_102_2_R0_data),
    .R0_en(mem_102_2_R0_en),
    .W0_addr(mem_102_2_W0_addr),
    .W0_clk(mem_102_2_W0_clk),
    .W0_data(mem_102_2_W0_data),
    .W0_en(mem_102_2_W0_en),
    .W0_mask(mem_102_2_W0_mask)
  );
  split_mem_0_ext mem_102_3 (
    .R0_addr(mem_102_3_R0_addr),
    .R0_clk(mem_102_3_R0_clk),
    .R0_data(mem_102_3_R0_data),
    .R0_en(mem_102_3_R0_en),
    .W0_addr(mem_102_3_W0_addr),
    .W0_clk(mem_102_3_W0_clk),
    .W0_data(mem_102_3_W0_data),
    .W0_en(mem_102_3_W0_en),
    .W0_mask(mem_102_3_W0_mask)
  );
  split_mem_0_ext mem_102_4 (
    .R0_addr(mem_102_4_R0_addr),
    .R0_clk(mem_102_4_R0_clk),
    .R0_data(mem_102_4_R0_data),
    .R0_en(mem_102_4_R0_en),
    .W0_addr(mem_102_4_W0_addr),
    .W0_clk(mem_102_4_W0_clk),
    .W0_data(mem_102_4_W0_data),
    .W0_en(mem_102_4_W0_en),
    .W0_mask(mem_102_4_W0_mask)
  );
  split_mem_0_ext mem_102_5 (
    .R0_addr(mem_102_5_R0_addr),
    .R0_clk(mem_102_5_R0_clk),
    .R0_data(mem_102_5_R0_data),
    .R0_en(mem_102_5_R0_en),
    .W0_addr(mem_102_5_W0_addr),
    .W0_clk(mem_102_5_W0_clk),
    .W0_data(mem_102_5_W0_data),
    .W0_en(mem_102_5_W0_en),
    .W0_mask(mem_102_5_W0_mask)
  );
  split_mem_0_ext mem_102_6 (
    .R0_addr(mem_102_6_R0_addr),
    .R0_clk(mem_102_6_R0_clk),
    .R0_data(mem_102_6_R0_data),
    .R0_en(mem_102_6_R0_en),
    .W0_addr(mem_102_6_W0_addr),
    .W0_clk(mem_102_6_W0_clk),
    .W0_data(mem_102_6_W0_data),
    .W0_en(mem_102_6_W0_en),
    .W0_mask(mem_102_6_W0_mask)
  );
  split_mem_0_ext mem_102_7 (
    .R0_addr(mem_102_7_R0_addr),
    .R0_clk(mem_102_7_R0_clk),
    .R0_data(mem_102_7_R0_data),
    .R0_en(mem_102_7_R0_en),
    .W0_addr(mem_102_7_W0_addr),
    .W0_clk(mem_102_7_W0_clk),
    .W0_data(mem_102_7_W0_data),
    .W0_en(mem_102_7_W0_en),
    .W0_mask(mem_102_7_W0_mask)
  );
  split_mem_0_ext mem_103_0 (
    .R0_addr(mem_103_0_R0_addr),
    .R0_clk(mem_103_0_R0_clk),
    .R0_data(mem_103_0_R0_data),
    .R0_en(mem_103_0_R0_en),
    .W0_addr(mem_103_0_W0_addr),
    .W0_clk(mem_103_0_W0_clk),
    .W0_data(mem_103_0_W0_data),
    .W0_en(mem_103_0_W0_en),
    .W0_mask(mem_103_0_W0_mask)
  );
  split_mem_0_ext mem_103_1 (
    .R0_addr(mem_103_1_R0_addr),
    .R0_clk(mem_103_1_R0_clk),
    .R0_data(mem_103_1_R0_data),
    .R0_en(mem_103_1_R0_en),
    .W0_addr(mem_103_1_W0_addr),
    .W0_clk(mem_103_1_W0_clk),
    .W0_data(mem_103_1_W0_data),
    .W0_en(mem_103_1_W0_en),
    .W0_mask(mem_103_1_W0_mask)
  );
  split_mem_0_ext mem_103_2 (
    .R0_addr(mem_103_2_R0_addr),
    .R0_clk(mem_103_2_R0_clk),
    .R0_data(mem_103_2_R0_data),
    .R0_en(mem_103_2_R0_en),
    .W0_addr(mem_103_2_W0_addr),
    .W0_clk(mem_103_2_W0_clk),
    .W0_data(mem_103_2_W0_data),
    .W0_en(mem_103_2_W0_en),
    .W0_mask(mem_103_2_W0_mask)
  );
  split_mem_0_ext mem_103_3 (
    .R0_addr(mem_103_3_R0_addr),
    .R0_clk(mem_103_3_R0_clk),
    .R0_data(mem_103_3_R0_data),
    .R0_en(mem_103_3_R0_en),
    .W0_addr(mem_103_3_W0_addr),
    .W0_clk(mem_103_3_W0_clk),
    .W0_data(mem_103_3_W0_data),
    .W0_en(mem_103_3_W0_en),
    .W0_mask(mem_103_3_W0_mask)
  );
  split_mem_0_ext mem_103_4 (
    .R0_addr(mem_103_4_R0_addr),
    .R0_clk(mem_103_4_R0_clk),
    .R0_data(mem_103_4_R0_data),
    .R0_en(mem_103_4_R0_en),
    .W0_addr(mem_103_4_W0_addr),
    .W0_clk(mem_103_4_W0_clk),
    .W0_data(mem_103_4_W0_data),
    .W0_en(mem_103_4_W0_en),
    .W0_mask(mem_103_4_W0_mask)
  );
  split_mem_0_ext mem_103_5 (
    .R0_addr(mem_103_5_R0_addr),
    .R0_clk(mem_103_5_R0_clk),
    .R0_data(mem_103_5_R0_data),
    .R0_en(mem_103_5_R0_en),
    .W0_addr(mem_103_5_W0_addr),
    .W0_clk(mem_103_5_W0_clk),
    .W0_data(mem_103_5_W0_data),
    .W0_en(mem_103_5_W0_en),
    .W0_mask(mem_103_5_W0_mask)
  );
  split_mem_0_ext mem_103_6 (
    .R0_addr(mem_103_6_R0_addr),
    .R0_clk(mem_103_6_R0_clk),
    .R0_data(mem_103_6_R0_data),
    .R0_en(mem_103_6_R0_en),
    .W0_addr(mem_103_6_W0_addr),
    .W0_clk(mem_103_6_W0_clk),
    .W0_data(mem_103_6_W0_data),
    .W0_en(mem_103_6_W0_en),
    .W0_mask(mem_103_6_W0_mask)
  );
  split_mem_0_ext mem_103_7 (
    .R0_addr(mem_103_7_R0_addr),
    .R0_clk(mem_103_7_R0_clk),
    .R0_data(mem_103_7_R0_data),
    .R0_en(mem_103_7_R0_en),
    .W0_addr(mem_103_7_W0_addr),
    .W0_clk(mem_103_7_W0_clk),
    .W0_data(mem_103_7_W0_data),
    .W0_en(mem_103_7_W0_en),
    .W0_mask(mem_103_7_W0_mask)
  );
  split_mem_0_ext mem_104_0 (
    .R0_addr(mem_104_0_R0_addr),
    .R0_clk(mem_104_0_R0_clk),
    .R0_data(mem_104_0_R0_data),
    .R0_en(mem_104_0_R0_en),
    .W0_addr(mem_104_0_W0_addr),
    .W0_clk(mem_104_0_W0_clk),
    .W0_data(mem_104_0_W0_data),
    .W0_en(mem_104_0_W0_en),
    .W0_mask(mem_104_0_W0_mask)
  );
  split_mem_0_ext mem_104_1 (
    .R0_addr(mem_104_1_R0_addr),
    .R0_clk(mem_104_1_R0_clk),
    .R0_data(mem_104_1_R0_data),
    .R0_en(mem_104_1_R0_en),
    .W0_addr(mem_104_1_W0_addr),
    .W0_clk(mem_104_1_W0_clk),
    .W0_data(mem_104_1_W0_data),
    .W0_en(mem_104_1_W0_en),
    .W0_mask(mem_104_1_W0_mask)
  );
  split_mem_0_ext mem_104_2 (
    .R0_addr(mem_104_2_R0_addr),
    .R0_clk(mem_104_2_R0_clk),
    .R0_data(mem_104_2_R0_data),
    .R0_en(mem_104_2_R0_en),
    .W0_addr(mem_104_2_W0_addr),
    .W0_clk(mem_104_2_W0_clk),
    .W0_data(mem_104_2_W0_data),
    .W0_en(mem_104_2_W0_en),
    .W0_mask(mem_104_2_W0_mask)
  );
  split_mem_0_ext mem_104_3 (
    .R0_addr(mem_104_3_R0_addr),
    .R0_clk(mem_104_3_R0_clk),
    .R0_data(mem_104_3_R0_data),
    .R0_en(mem_104_3_R0_en),
    .W0_addr(mem_104_3_W0_addr),
    .W0_clk(mem_104_3_W0_clk),
    .W0_data(mem_104_3_W0_data),
    .W0_en(mem_104_3_W0_en),
    .W0_mask(mem_104_3_W0_mask)
  );
  split_mem_0_ext mem_104_4 (
    .R0_addr(mem_104_4_R0_addr),
    .R0_clk(mem_104_4_R0_clk),
    .R0_data(mem_104_4_R0_data),
    .R0_en(mem_104_4_R0_en),
    .W0_addr(mem_104_4_W0_addr),
    .W0_clk(mem_104_4_W0_clk),
    .W0_data(mem_104_4_W0_data),
    .W0_en(mem_104_4_W0_en),
    .W0_mask(mem_104_4_W0_mask)
  );
  split_mem_0_ext mem_104_5 (
    .R0_addr(mem_104_5_R0_addr),
    .R0_clk(mem_104_5_R0_clk),
    .R0_data(mem_104_5_R0_data),
    .R0_en(mem_104_5_R0_en),
    .W0_addr(mem_104_5_W0_addr),
    .W0_clk(mem_104_5_W0_clk),
    .W0_data(mem_104_5_W0_data),
    .W0_en(mem_104_5_W0_en),
    .W0_mask(mem_104_5_W0_mask)
  );
  split_mem_0_ext mem_104_6 (
    .R0_addr(mem_104_6_R0_addr),
    .R0_clk(mem_104_6_R0_clk),
    .R0_data(mem_104_6_R0_data),
    .R0_en(mem_104_6_R0_en),
    .W0_addr(mem_104_6_W0_addr),
    .W0_clk(mem_104_6_W0_clk),
    .W0_data(mem_104_6_W0_data),
    .W0_en(mem_104_6_W0_en),
    .W0_mask(mem_104_6_W0_mask)
  );
  split_mem_0_ext mem_104_7 (
    .R0_addr(mem_104_7_R0_addr),
    .R0_clk(mem_104_7_R0_clk),
    .R0_data(mem_104_7_R0_data),
    .R0_en(mem_104_7_R0_en),
    .W0_addr(mem_104_7_W0_addr),
    .W0_clk(mem_104_7_W0_clk),
    .W0_data(mem_104_7_W0_data),
    .W0_en(mem_104_7_W0_en),
    .W0_mask(mem_104_7_W0_mask)
  );
  split_mem_0_ext mem_105_0 (
    .R0_addr(mem_105_0_R0_addr),
    .R0_clk(mem_105_0_R0_clk),
    .R0_data(mem_105_0_R0_data),
    .R0_en(mem_105_0_R0_en),
    .W0_addr(mem_105_0_W0_addr),
    .W0_clk(mem_105_0_W0_clk),
    .W0_data(mem_105_0_W0_data),
    .W0_en(mem_105_0_W0_en),
    .W0_mask(mem_105_0_W0_mask)
  );
  split_mem_0_ext mem_105_1 (
    .R0_addr(mem_105_1_R0_addr),
    .R0_clk(mem_105_1_R0_clk),
    .R0_data(mem_105_1_R0_data),
    .R0_en(mem_105_1_R0_en),
    .W0_addr(mem_105_1_W0_addr),
    .W0_clk(mem_105_1_W0_clk),
    .W0_data(mem_105_1_W0_data),
    .W0_en(mem_105_1_W0_en),
    .W0_mask(mem_105_1_W0_mask)
  );
  split_mem_0_ext mem_105_2 (
    .R0_addr(mem_105_2_R0_addr),
    .R0_clk(mem_105_2_R0_clk),
    .R0_data(mem_105_2_R0_data),
    .R0_en(mem_105_2_R0_en),
    .W0_addr(mem_105_2_W0_addr),
    .W0_clk(mem_105_2_W0_clk),
    .W0_data(mem_105_2_W0_data),
    .W0_en(mem_105_2_W0_en),
    .W0_mask(mem_105_2_W0_mask)
  );
  split_mem_0_ext mem_105_3 (
    .R0_addr(mem_105_3_R0_addr),
    .R0_clk(mem_105_3_R0_clk),
    .R0_data(mem_105_3_R0_data),
    .R0_en(mem_105_3_R0_en),
    .W0_addr(mem_105_3_W0_addr),
    .W0_clk(mem_105_3_W0_clk),
    .W0_data(mem_105_3_W0_data),
    .W0_en(mem_105_3_W0_en),
    .W0_mask(mem_105_3_W0_mask)
  );
  split_mem_0_ext mem_105_4 (
    .R0_addr(mem_105_4_R0_addr),
    .R0_clk(mem_105_4_R0_clk),
    .R0_data(mem_105_4_R0_data),
    .R0_en(mem_105_4_R0_en),
    .W0_addr(mem_105_4_W0_addr),
    .W0_clk(mem_105_4_W0_clk),
    .W0_data(mem_105_4_W0_data),
    .W0_en(mem_105_4_W0_en),
    .W0_mask(mem_105_4_W0_mask)
  );
  split_mem_0_ext mem_105_5 (
    .R0_addr(mem_105_5_R0_addr),
    .R0_clk(mem_105_5_R0_clk),
    .R0_data(mem_105_5_R0_data),
    .R0_en(mem_105_5_R0_en),
    .W0_addr(mem_105_5_W0_addr),
    .W0_clk(mem_105_5_W0_clk),
    .W0_data(mem_105_5_W0_data),
    .W0_en(mem_105_5_W0_en),
    .W0_mask(mem_105_5_W0_mask)
  );
  split_mem_0_ext mem_105_6 (
    .R0_addr(mem_105_6_R0_addr),
    .R0_clk(mem_105_6_R0_clk),
    .R0_data(mem_105_6_R0_data),
    .R0_en(mem_105_6_R0_en),
    .W0_addr(mem_105_6_W0_addr),
    .W0_clk(mem_105_6_W0_clk),
    .W0_data(mem_105_6_W0_data),
    .W0_en(mem_105_6_W0_en),
    .W0_mask(mem_105_6_W0_mask)
  );
  split_mem_0_ext mem_105_7 (
    .R0_addr(mem_105_7_R0_addr),
    .R0_clk(mem_105_7_R0_clk),
    .R0_data(mem_105_7_R0_data),
    .R0_en(mem_105_7_R0_en),
    .W0_addr(mem_105_7_W0_addr),
    .W0_clk(mem_105_7_W0_clk),
    .W0_data(mem_105_7_W0_data),
    .W0_en(mem_105_7_W0_en),
    .W0_mask(mem_105_7_W0_mask)
  );
  split_mem_0_ext mem_106_0 (
    .R0_addr(mem_106_0_R0_addr),
    .R0_clk(mem_106_0_R0_clk),
    .R0_data(mem_106_0_R0_data),
    .R0_en(mem_106_0_R0_en),
    .W0_addr(mem_106_0_W0_addr),
    .W0_clk(mem_106_0_W0_clk),
    .W0_data(mem_106_0_W0_data),
    .W0_en(mem_106_0_W0_en),
    .W0_mask(mem_106_0_W0_mask)
  );
  split_mem_0_ext mem_106_1 (
    .R0_addr(mem_106_1_R0_addr),
    .R0_clk(mem_106_1_R0_clk),
    .R0_data(mem_106_1_R0_data),
    .R0_en(mem_106_1_R0_en),
    .W0_addr(mem_106_1_W0_addr),
    .W0_clk(mem_106_1_W0_clk),
    .W0_data(mem_106_1_W0_data),
    .W0_en(mem_106_1_W0_en),
    .W0_mask(mem_106_1_W0_mask)
  );
  split_mem_0_ext mem_106_2 (
    .R0_addr(mem_106_2_R0_addr),
    .R0_clk(mem_106_2_R0_clk),
    .R0_data(mem_106_2_R0_data),
    .R0_en(mem_106_2_R0_en),
    .W0_addr(mem_106_2_W0_addr),
    .W0_clk(mem_106_2_W0_clk),
    .W0_data(mem_106_2_W0_data),
    .W0_en(mem_106_2_W0_en),
    .W0_mask(mem_106_2_W0_mask)
  );
  split_mem_0_ext mem_106_3 (
    .R0_addr(mem_106_3_R0_addr),
    .R0_clk(mem_106_3_R0_clk),
    .R0_data(mem_106_3_R0_data),
    .R0_en(mem_106_3_R0_en),
    .W0_addr(mem_106_3_W0_addr),
    .W0_clk(mem_106_3_W0_clk),
    .W0_data(mem_106_3_W0_data),
    .W0_en(mem_106_3_W0_en),
    .W0_mask(mem_106_3_W0_mask)
  );
  split_mem_0_ext mem_106_4 (
    .R0_addr(mem_106_4_R0_addr),
    .R0_clk(mem_106_4_R0_clk),
    .R0_data(mem_106_4_R0_data),
    .R0_en(mem_106_4_R0_en),
    .W0_addr(mem_106_4_W0_addr),
    .W0_clk(mem_106_4_W0_clk),
    .W0_data(mem_106_4_W0_data),
    .W0_en(mem_106_4_W0_en),
    .W0_mask(mem_106_4_W0_mask)
  );
  split_mem_0_ext mem_106_5 (
    .R0_addr(mem_106_5_R0_addr),
    .R0_clk(mem_106_5_R0_clk),
    .R0_data(mem_106_5_R0_data),
    .R0_en(mem_106_5_R0_en),
    .W0_addr(mem_106_5_W0_addr),
    .W0_clk(mem_106_5_W0_clk),
    .W0_data(mem_106_5_W0_data),
    .W0_en(mem_106_5_W0_en),
    .W0_mask(mem_106_5_W0_mask)
  );
  split_mem_0_ext mem_106_6 (
    .R0_addr(mem_106_6_R0_addr),
    .R0_clk(mem_106_6_R0_clk),
    .R0_data(mem_106_6_R0_data),
    .R0_en(mem_106_6_R0_en),
    .W0_addr(mem_106_6_W0_addr),
    .W0_clk(mem_106_6_W0_clk),
    .W0_data(mem_106_6_W0_data),
    .W0_en(mem_106_6_W0_en),
    .W0_mask(mem_106_6_W0_mask)
  );
  split_mem_0_ext mem_106_7 (
    .R0_addr(mem_106_7_R0_addr),
    .R0_clk(mem_106_7_R0_clk),
    .R0_data(mem_106_7_R0_data),
    .R0_en(mem_106_7_R0_en),
    .W0_addr(mem_106_7_W0_addr),
    .W0_clk(mem_106_7_W0_clk),
    .W0_data(mem_106_7_W0_data),
    .W0_en(mem_106_7_W0_en),
    .W0_mask(mem_106_7_W0_mask)
  );
  split_mem_0_ext mem_107_0 (
    .R0_addr(mem_107_0_R0_addr),
    .R0_clk(mem_107_0_R0_clk),
    .R0_data(mem_107_0_R0_data),
    .R0_en(mem_107_0_R0_en),
    .W0_addr(mem_107_0_W0_addr),
    .W0_clk(mem_107_0_W0_clk),
    .W0_data(mem_107_0_W0_data),
    .W0_en(mem_107_0_W0_en),
    .W0_mask(mem_107_0_W0_mask)
  );
  split_mem_0_ext mem_107_1 (
    .R0_addr(mem_107_1_R0_addr),
    .R0_clk(mem_107_1_R0_clk),
    .R0_data(mem_107_1_R0_data),
    .R0_en(mem_107_1_R0_en),
    .W0_addr(mem_107_1_W0_addr),
    .W0_clk(mem_107_1_W0_clk),
    .W0_data(mem_107_1_W0_data),
    .W0_en(mem_107_1_W0_en),
    .W0_mask(mem_107_1_W0_mask)
  );
  split_mem_0_ext mem_107_2 (
    .R0_addr(mem_107_2_R0_addr),
    .R0_clk(mem_107_2_R0_clk),
    .R0_data(mem_107_2_R0_data),
    .R0_en(mem_107_2_R0_en),
    .W0_addr(mem_107_2_W0_addr),
    .W0_clk(mem_107_2_W0_clk),
    .W0_data(mem_107_2_W0_data),
    .W0_en(mem_107_2_W0_en),
    .W0_mask(mem_107_2_W0_mask)
  );
  split_mem_0_ext mem_107_3 (
    .R0_addr(mem_107_3_R0_addr),
    .R0_clk(mem_107_3_R0_clk),
    .R0_data(mem_107_3_R0_data),
    .R0_en(mem_107_3_R0_en),
    .W0_addr(mem_107_3_W0_addr),
    .W0_clk(mem_107_3_W0_clk),
    .W0_data(mem_107_3_W0_data),
    .W0_en(mem_107_3_W0_en),
    .W0_mask(mem_107_3_W0_mask)
  );
  split_mem_0_ext mem_107_4 (
    .R0_addr(mem_107_4_R0_addr),
    .R0_clk(mem_107_4_R0_clk),
    .R0_data(mem_107_4_R0_data),
    .R0_en(mem_107_4_R0_en),
    .W0_addr(mem_107_4_W0_addr),
    .W0_clk(mem_107_4_W0_clk),
    .W0_data(mem_107_4_W0_data),
    .W0_en(mem_107_4_W0_en),
    .W0_mask(mem_107_4_W0_mask)
  );
  split_mem_0_ext mem_107_5 (
    .R0_addr(mem_107_5_R0_addr),
    .R0_clk(mem_107_5_R0_clk),
    .R0_data(mem_107_5_R0_data),
    .R0_en(mem_107_5_R0_en),
    .W0_addr(mem_107_5_W0_addr),
    .W0_clk(mem_107_5_W0_clk),
    .W0_data(mem_107_5_W0_data),
    .W0_en(mem_107_5_W0_en),
    .W0_mask(mem_107_5_W0_mask)
  );
  split_mem_0_ext mem_107_6 (
    .R0_addr(mem_107_6_R0_addr),
    .R0_clk(mem_107_6_R0_clk),
    .R0_data(mem_107_6_R0_data),
    .R0_en(mem_107_6_R0_en),
    .W0_addr(mem_107_6_W0_addr),
    .W0_clk(mem_107_6_W0_clk),
    .W0_data(mem_107_6_W0_data),
    .W0_en(mem_107_6_W0_en),
    .W0_mask(mem_107_6_W0_mask)
  );
  split_mem_0_ext mem_107_7 (
    .R0_addr(mem_107_7_R0_addr),
    .R0_clk(mem_107_7_R0_clk),
    .R0_data(mem_107_7_R0_data),
    .R0_en(mem_107_7_R0_en),
    .W0_addr(mem_107_7_W0_addr),
    .W0_clk(mem_107_7_W0_clk),
    .W0_data(mem_107_7_W0_data),
    .W0_en(mem_107_7_W0_en),
    .W0_mask(mem_107_7_W0_mask)
  );
  split_mem_0_ext mem_108_0 (
    .R0_addr(mem_108_0_R0_addr),
    .R0_clk(mem_108_0_R0_clk),
    .R0_data(mem_108_0_R0_data),
    .R0_en(mem_108_0_R0_en),
    .W0_addr(mem_108_0_W0_addr),
    .W0_clk(mem_108_0_W0_clk),
    .W0_data(mem_108_0_W0_data),
    .W0_en(mem_108_0_W0_en),
    .W0_mask(mem_108_0_W0_mask)
  );
  split_mem_0_ext mem_108_1 (
    .R0_addr(mem_108_1_R0_addr),
    .R0_clk(mem_108_1_R0_clk),
    .R0_data(mem_108_1_R0_data),
    .R0_en(mem_108_1_R0_en),
    .W0_addr(mem_108_1_W0_addr),
    .W0_clk(mem_108_1_W0_clk),
    .W0_data(mem_108_1_W0_data),
    .W0_en(mem_108_1_W0_en),
    .W0_mask(mem_108_1_W0_mask)
  );
  split_mem_0_ext mem_108_2 (
    .R0_addr(mem_108_2_R0_addr),
    .R0_clk(mem_108_2_R0_clk),
    .R0_data(mem_108_2_R0_data),
    .R0_en(mem_108_2_R0_en),
    .W0_addr(mem_108_2_W0_addr),
    .W0_clk(mem_108_2_W0_clk),
    .W0_data(mem_108_2_W0_data),
    .W0_en(mem_108_2_W0_en),
    .W0_mask(mem_108_2_W0_mask)
  );
  split_mem_0_ext mem_108_3 (
    .R0_addr(mem_108_3_R0_addr),
    .R0_clk(mem_108_3_R0_clk),
    .R0_data(mem_108_3_R0_data),
    .R0_en(mem_108_3_R0_en),
    .W0_addr(mem_108_3_W0_addr),
    .W0_clk(mem_108_3_W0_clk),
    .W0_data(mem_108_3_W0_data),
    .W0_en(mem_108_3_W0_en),
    .W0_mask(mem_108_3_W0_mask)
  );
  split_mem_0_ext mem_108_4 (
    .R0_addr(mem_108_4_R0_addr),
    .R0_clk(mem_108_4_R0_clk),
    .R0_data(mem_108_4_R0_data),
    .R0_en(mem_108_4_R0_en),
    .W0_addr(mem_108_4_W0_addr),
    .W0_clk(mem_108_4_W0_clk),
    .W0_data(mem_108_4_W0_data),
    .W0_en(mem_108_4_W0_en),
    .W0_mask(mem_108_4_W0_mask)
  );
  split_mem_0_ext mem_108_5 (
    .R0_addr(mem_108_5_R0_addr),
    .R0_clk(mem_108_5_R0_clk),
    .R0_data(mem_108_5_R0_data),
    .R0_en(mem_108_5_R0_en),
    .W0_addr(mem_108_5_W0_addr),
    .W0_clk(mem_108_5_W0_clk),
    .W0_data(mem_108_5_W0_data),
    .W0_en(mem_108_5_W0_en),
    .W0_mask(mem_108_5_W0_mask)
  );
  split_mem_0_ext mem_108_6 (
    .R0_addr(mem_108_6_R0_addr),
    .R0_clk(mem_108_6_R0_clk),
    .R0_data(mem_108_6_R0_data),
    .R0_en(mem_108_6_R0_en),
    .W0_addr(mem_108_6_W0_addr),
    .W0_clk(mem_108_6_W0_clk),
    .W0_data(mem_108_6_W0_data),
    .W0_en(mem_108_6_W0_en),
    .W0_mask(mem_108_6_W0_mask)
  );
  split_mem_0_ext mem_108_7 (
    .R0_addr(mem_108_7_R0_addr),
    .R0_clk(mem_108_7_R0_clk),
    .R0_data(mem_108_7_R0_data),
    .R0_en(mem_108_7_R0_en),
    .W0_addr(mem_108_7_W0_addr),
    .W0_clk(mem_108_7_W0_clk),
    .W0_data(mem_108_7_W0_data),
    .W0_en(mem_108_7_W0_en),
    .W0_mask(mem_108_7_W0_mask)
  );
  split_mem_0_ext mem_109_0 (
    .R0_addr(mem_109_0_R0_addr),
    .R0_clk(mem_109_0_R0_clk),
    .R0_data(mem_109_0_R0_data),
    .R0_en(mem_109_0_R0_en),
    .W0_addr(mem_109_0_W0_addr),
    .W0_clk(mem_109_0_W0_clk),
    .W0_data(mem_109_0_W0_data),
    .W0_en(mem_109_0_W0_en),
    .W0_mask(mem_109_0_W0_mask)
  );
  split_mem_0_ext mem_109_1 (
    .R0_addr(mem_109_1_R0_addr),
    .R0_clk(mem_109_1_R0_clk),
    .R0_data(mem_109_1_R0_data),
    .R0_en(mem_109_1_R0_en),
    .W0_addr(mem_109_1_W0_addr),
    .W0_clk(mem_109_1_W0_clk),
    .W0_data(mem_109_1_W0_data),
    .W0_en(mem_109_1_W0_en),
    .W0_mask(mem_109_1_W0_mask)
  );
  split_mem_0_ext mem_109_2 (
    .R0_addr(mem_109_2_R0_addr),
    .R0_clk(mem_109_2_R0_clk),
    .R0_data(mem_109_2_R0_data),
    .R0_en(mem_109_2_R0_en),
    .W0_addr(mem_109_2_W0_addr),
    .W0_clk(mem_109_2_W0_clk),
    .W0_data(mem_109_2_W0_data),
    .W0_en(mem_109_2_W0_en),
    .W0_mask(mem_109_2_W0_mask)
  );
  split_mem_0_ext mem_109_3 (
    .R0_addr(mem_109_3_R0_addr),
    .R0_clk(mem_109_3_R0_clk),
    .R0_data(mem_109_3_R0_data),
    .R0_en(mem_109_3_R0_en),
    .W0_addr(mem_109_3_W0_addr),
    .W0_clk(mem_109_3_W0_clk),
    .W0_data(mem_109_3_W0_data),
    .W0_en(mem_109_3_W0_en),
    .W0_mask(mem_109_3_W0_mask)
  );
  split_mem_0_ext mem_109_4 (
    .R0_addr(mem_109_4_R0_addr),
    .R0_clk(mem_109_4_R0_clk),
    .R0_data(mem_109_4_R0_data),
    .R0_en(mem_109_4_R0_en),
    .W0_addr(mem_109_4_W0_addr),
    .W0_clk(mem_109_4_W0_clk),
    .W0_data(mem_109_4_W0_data),
    .W0_en(mem_109_4_W0_en),
    .W0_mask(mem_109_4_W0_mask)
  );
  split_mem_0_ext mem_109_5 (
    .R0_addr(mem_109_5_R0_addr),
    .R0_clk(mem_109_5_R0_clk),
    .R0_data(mem_109_5_R0_data),
    .R0_en(mem_109_5_R0_en),
    .W0_addr(mem_109_5_W0_addr),
    .W0_clk(mem_109_5_W0_clk),
    .W0_data(mem_109_5_W0_data),
    .W0_en(mem_109_5_W0_en),
    .W0_mask(mem_109_5_W0_mask)
  );
  split_mem_0_ext mem_109_6 (
    .R0_addr(mem_109_6_R0_addr),
    .R0_clk(mem_109_6_R0_clk),
    .R0_data(mem_109_6_R0_data),
    .R0_en(mem_109_6_R0_en),
    .W0_addr(mem_109_6_W0_addr),
    .W0_clk(mem_109_6_W0_clk),
    .W0_data(mem_109_6_W0_data),
    .W0_en(mem_109_6_W0_en),
    .W0_mask(mem_109_6_W0_mask)
  );
  split_mem_0_ext mem_109_7 (
    .R0_addr(mem_109_7_R0_addr),
    .R0_clk(mem_109_7_R0_clk),
    .R0_data(mem_109_7_R0_data),
    .R0_en(mem_109_7_R0_en),
    .W0_addr(mem_109_7_W0_addr),
    .W0_clk(mem_109_7_W0_clk),
    .W0_data(mem_109_7_W0_data),
    .W0_en(mem_109_7_W0_en),
    .W0_mask(mem_109_7_W0_mask)
  );
  split_mem_0_ext mem_110_0 (
    .R0_addr(mem_110_0_R0_addr),
    .R0_clk(mem_110_0_R0_clk),
    .R0_data(mem_110_0_R0_data),
    .R0_en(mem_110_0_R0_en),
    .W0_addr(mem_110_0_W0_addr),
    .W0_clk(mem_110_0_W0_clk),
    .W0_data(mem_110_0_W0_data),
    .W0_en(mem_110_0_W0_en),
    .W0_mask(mem_110_0_W0_mask)
  );
  split_mem_0_ext mem_110_1 (
    .R0_addr(mem_110_1_R0_addr),
    .R0_clk(mem_110_1_R0_clk),
    .R0_data(mem_110_1_R0_data),
    .R0_en(mem_110_1_R0_en),
    .W0_addr(mem_110_1_W0_addr),
    .W0_clk(mem_110_1_W0_clk),
    .W0_data(mem_110_1_W0_data),
    .W0_en(mem_110_1_W0_en),
    .W0_mask(mem_110_1_W0_mask)
  );
  split_mem_0_ext mem_110_2 (
    .R0_addr(mem_110_2_R0_addr),
    .R0_clk(mem_110_2_R0_clk),
    .R0_data(mem_110_2_R0_data),
    .R0_en(mem_110_2_R0_en),
    .W0_addr(mem_110_2_W0_addr),
    .W0_clk(mem_110_2_W0_clk),
    .W0_data(mem_110_2_W0_data),
    .W0_en(mem_110_2_W0_en),
    .W0_mask(mem_110_2_W0_mask)
  );
  split_mem_0_ext mem_110_3 (
    .R0_addr(mem_110_3_R0_addr),
    .R0_clk(mem_110_3_R0_clk),
    .R0_data(mem_110_3_R0_data),
    .R0_en(mem_110_3_R0_en),
    .W0_addr(mem_110_3_W0_addr),
    .W0_clk(mem_110_3_W0_clk),
    .W0_data(mem_110_3_W0_data),
    .W0_en(mem_110_3_W0_en),
    .W0_mask(mem_110_3_W0_mask)
  );
  split_mem_0_ext mem_110_4 (
    .R0_addr(mem_110_4_R0_addr),
    .R0_clk(mem_110_4_R0_clk),
    .R0_data(mem_110_4_R0_data),
    .R0_en(mem_110_4_R0_en),
    .W0_addr(mem_110_4_W0_addr),
    .W0_clk(mem_110_4_W0_clk),
    .W0_data(mem_110_4_W0_data),
    .W0_en(mem_110_4_W0_en),
    .W0_mask(mem_110_4_W0_mask)
  );
  split_mem_0_ext mem_110_5 (
    .R0_addr(mem_110_5_R0_addr),
    .R0_clk(mem_110_5_R0_clk),
    .R0_data(mem_110_5_R0_data),
    .R0_en(mem_110_5_R0_en),
    .W0_addr(mem_110_5_W0_addr),
    .W0_clk(mem_110_5_W0_clk),
    .W0_data(mem_110_5_W0_data),
    .W0_en(mem_110_5_W0_en),
    .W0_mask(mem_110_5_W0_mask)
  );
  split_mem_0_ext mem_110_6 (
    .R0_addr(mem_110_6_R0_addr),
    .R0_clk(mem_110_6_R0_clk),
    .R0_data(mem_110_6_R0_data),
    .R0_en(mem_110_6_R0_en),
    .W0_addr(mem_110_6_W0_addr),
    .W0_clk(mem_110_6_W0_clk),
    .W0_data(mem_110_6_W0_data),
    .W0_en(mem_110_6_W0_en),
    .W0_mask(mem_110_6_W0_mask)
  );
  split_mem_0_ext mem_110_7 (
    .R0_addr(mem_110_7_R0_addr),
    .R0_clk(mem_110_7_R0_clk),
    .R0_data(mem_110_7_R0_data),
    .R0_en(mem_110_7_R0_en),
    .W0_addr(mem_110_7_W0_addr),
    .W0_clk(mem_110_7_W0_clk),
    .W0_data(mem_110_7_W0_data),
    .W0_en(mem_110_7_W0_en),
    .W0_mask(mem_110_7_W0_mask)
  );
  split_mem_0_ext mem_111_0 (
    .R0_addr(mem_111_0_R0_addr),
    .R0_clk(mem_111_0_R0_clk),
    .R0_data(mem_111_0_R0_data),
    .R0_en(mem_111_0_R0_en),
    .W0_addr(mem_111_0_W0_addr),
    .W0_clk(mem_111_0_W0_clk),
    .W0_data(mem_111_0_W0_data),
    .W0_en(mem_111_0_W0_en),
    .W0_mask(mem_111_0_W0_mask)
  );
  split_mem_0_ext mem_111_1 (
    .R0_addr(mem_111_1_R0_addr),
    .R0_clk(mem_111_1_R0_clk),
    .R0_data(mem_111_1_R0_data),
    .R0_en(mem_111_1_R0_en),
    .W0_addr(mem_111_1_W0_addr),
    .W0_clk(mem_111_1_W0_clk),
    .W0_data(mem_111_1_W0_data),
    .W0_en(mem_111_1_W0_en),
    .W0_mask(mem_111_1_W0_mask)
  );
  split_mem_0_ext mem_111_2 (
    .R0_addr(mem_111_2_R0_addr),
    .R0_clk(mem_111_2_R0_clk),
    .R0_data(mem_111_2_R0_data),
    .R0_en(mem_111_2_R0_en),
    .W0_addr(mem_111_2_W0_addr),
    .W0_clk(mem_111_2_W0_clk),
    .W0_data(mem_111_2_W0_data),
    .W0_en(mem_111_2_W0_en),
    .W0_mask(mem_111_2_W0_mask)
  );
  split_mem_0_ext mem_111_3 (
    .R0_addr(mem_111_3_R0_addr),
    .R0_clk(mem_111_3_R0_clk),
    .R0_data(mem_111_3_R0_data),
    .R0_en(mem_111_3_R0_en),
    .W0_addr(mem_111_3_W0_addr),
    .W0_clk(mem_111_3_W0_clk),
    .W0_data(mem_111_3_W0_data),
    .W0_en(mem_111_3_W0_en),
    .W0_mask(mem_111_3_W0_mask)
  );
  split_mem_0_ext mem_111_4 (
    .R0_addr(mem_111_4_R0_addr),
    .R0_clk(mem_111_4_R0_clk),
    .R0_data(mem_111_4_R0_data),
    .R0_en(mem_111_4_R0_en),
    .W0_addr(mem_111_4_W0_addr),
    .W0_clk(mem_111_4_W0_clk),
    .W0_data(mem_111_4_W0_data),
    .W0_en(mem_111_4_W0_en),
    .W0_mask(mem_111_4_W0_mask)
  );
  split_mem_0_ext mem_111_5 (
    .R0_addr(mem_111_5_R0_addr),
    .R0_clk(mem_111_5_R0_clk),
    .R0_data(mem_111_5_R0_data),
    .R0_en(mem_111_5_R0_en),
    .W0_addr(mem_111_5_W0_addr),
    .W0_clk(mem_111_5_W0_clk),
    .W0_data(mem_111_5_W0_data),
    .W0_en(mem_111_5_W0_en),
    .W0_mask(mem_111_5_W0_mask)
  );
  split_mem_0_ext mem_111_6 (
    .R0_addr(mem_111_6_R0_addr),
    .R0_clk(mem_111_6_R0_clk),
    .R0_data(mem_111_6_R0_data),
    .R0_en(mem_111_6_R0_en),
    .W0_addr(mem_111_6_W0_addr),
    .W0_clk(mem_111_6_W0_clk),
    .W0_data(mem_111_6_W0_data),
    .W0_en(mem_111_6_W0_en),
    .W0_mask(mem_111_6_W0_mask)
  );
  split_mem_0_ext mem_111_7 (
    .R0_addr(mem_111_7_R0_addr),
    .R0_clk(mem_111_7_R0_clk),
    .R0_data(mem_111_7_R0_data),
    .R0_en(mem_111_7_R0_en),
    .W0_addr(mem_111_7_W0_addr),
    .W0_clk(mem_111_7_W0_clk),
    .W0_data(mem_111_7_W0_data),
    .W0_en(mem_111_7_W0_en),
    .W0_mask(mem_111_7_W0_mask)
  );
  split_mem_0_ext mem_112_0 (
    .R0_addr(mem_112_0_R0_addr),
    .R0_clk(mem_112_0_R0_clk),
    .R0_data(mem_112_0_R0_data),
    .R0_en(mem_112_0_R0_en),
    .W0_addr(mem_112_0_W0_addr),
    .W0_clk(mem_112_0_W0_clk),
    .W0_data(mem_112_0_W0_data),
    .W0_en(mem_112_0_W0_en),
    .W0_mask(mem_112_0_W0_mask)
  );
  split_mem_0_ext mem_112_1 (
    .R0_addr(mem_112_1_R0_addr),
    .R0_clk(mem_112_1_R0_clk),
    .R0_data(mem_112_1_R0_data),
    .R0_en(mem_112_1_R0_en),
    .W0_addr(mem_112_1_W0_addr),
    .W0_clk(mem_112_1_W0_clk),
    .W0_data(mem_112_1_W0_data),
    .W0_en(mem_112_1_W0_en),
    .W0_mask(mem_112_1_W0_mask)
  );
  split_mem_0_ext mem_112_2 (
    .R0_addr(mem_112_2_R0_addr),
    .R0_clk(mem_112_2_R0_clk),
    .R0_data(mem_112_2_R0_data),
    .R0_en(mem_112_2_R0_en),
    .W0_addr(mem_112_2_W0_addr),
    .W0_clk(mem_112_2_W0_clk),
    .W0_data(mem_112_2_W0_data),
    .W0_en(mem_112_2_W0_en),
    .W0_mask(mem_112_2_W0_mask)
  );
  split_mem_0_ext mem_112_3 (
    .R0_addr(mem_112_3_R0_addr),
    .R0_clk(mem_112_3_R0_clk),
    .R0_data(mem_112_3_R0_data),
    .R0_en(mem_112_3_R0_en),
    .W0_addr(mem_112_3_W0_addr),
    .W0_clk(mem_112_3_W0_clk),
    .W0_data(mem_112_3_W0_data),
    .W0_en(mem_112_3_W0_en),
    .W0_mask(mem_112_3_W0_mask)
  );
  split_mem_0_ext mem_112_4 (
    .R0_addr(mem_112_4_R0_addr),
    .R0_clk(mem_112_4_R0_clk),
    .R0_data(mem_112_4_R0_data),
    .R0_en(mem_112_4_R0_en),
    .W0_addr(mem_112_4_W0_addr),
    .W0_clk(mem_112_4_W0_clk),
    .W0_data(mem_112_4_W0_data),
    .W0_en(mem_112_4_W0_en),
    .W0_mask(mem_112_4_W0_mask)
  );
  split_mem_0_ext mem_112_5 (
    .R0_addr(mem_112_5_R0_addr),
    .R0_clk(mem_112_5_R0_clk),
    .R0_data(mem_112_5_R0_data),
    .R0_en(mem_112_5_R0_en),
    .W0_addr(mem_112_5_W0_addr),
    .W0_clk(mem_112_5_W0_clk),
    .W0_data(mem_112_5_W0_data),
    .W0_en(mem_112_5_W0_en),
    .W0_mask(mem_112_5_W0_mask)
  );
  split_mem_0_ext mem_112_6 (
    .R0_addr(mem_112_6_R0_addr),
    .R0_clk(mem_112_6_R0_clk),
    .R0_data(mem_112_6_R0_data),
    .R0_en(mem_112_6_R0_en),
    .W0_addr(mem_112_6_W0_addr),
    .W0_clk(mem_112_6_W0_clk),
    .W0_data(mem_112_6_W0_data),
    .W0_en(mem_112_6_W0_en),
    .W0_mask(mem_112_6_W0_mask)
  );
  split_mem_0_ext mem_112_7 (
    .R0_addr(mem_112_7_R0_addr),
    .R0_clk(mem_112_7_R0_clk),
    .R0_data(mem_112_7_R0_data),
    .R0_en(mem_112_7_R0_en),
    .W0_addr(mem_112_7_W0_addr),
    .W0_clk(mem_112_7_W0_clk),
    .W0_data(mem_112_7_W0_data),
    .W0_en(mem_112_7_W0_en),
    .W0_mask(mem_112_7_W0_mask)
  );
  split_mem_0_ext mem_113_0 (
    .R0_addr(mem_113_0_R0_addr),
    .R0_clk(mem_113_0_R0_clk),
    .R0_data(mem_113_0_R0_data),
    .R0_en(mem_113_0_R0_en),
    .W0_addr(mem_113_0_W0_addr),
    .W0_clk(mem_113_0_W0_clk),
    .W0_data(mem_113_0_W0_data),
    .W0_en(mem_113_0_W0_en),
    .W0_mask(mem_113_0_W0_mask)
  );
  split_mem_0_ext mem_113_1 (
    .R0_addr(mem_113_1_R0_addr),
    .R0_clk(mem_113_1_R0_clk),
    .R0_data(mem_113_1_R0_data),
    .R0_en(mem_113_1_R0_en),
    .W0_addr(mem_113_1_W0_addr),
    .W0_clk(mem_113_1_W0_clk),
    .W0_data(mem_113_1_W0_data),
    .W0_en(mem_113_1_W0_en),
    .W0_mask(mem_113_1_W0_mask)
  );
  split_mem_0_ext mem_113_2 (
    .R0_addr(mem_113_2_R0_addr),
    .R0_clk(mem_113_2_R0_clk),
    .R0_data(mem_113_2_R0_data),
    .R0_en(mem_113_2_R0_en),
    .W0_addr(mem_113_2_W0_addr),
    .W0_clk(mem_113_2_W0_clk),
    .W0_data(mem_113_2_W0_data),
    .W0_en(mem_113_2_W0_en),
    .W0_mask(mem_113_2_W0_mask)
  );
  split_mem_0_ext mem_113_3 (
    .R0_addr(mem_113_3_R0_addr),
    .R0_clk(mem_113_3_R0_clk),
    .R0_data(mem_113_3_R0_data),
    .R0_en(mem_113_3_R0_en),
    .W0_addr(mem_113_3_W0_addr),
    .W0_clk(mem_113_3_W0_clk),
    .W0_data(mem_113_3_W0_data),
    .W0_en(mem_113_3_W0_en),
    .W0_mask(mem_113_3_W0_mask)
  );
  split_mem_0_ext mem_113_4 (
    .R0_addr(mem_113_4_R0_addr),
    .R0_clk(mem_113_4_R0_clk),
    .R0_data(mem_113_4_R0_data),
    .R0_en(mem_113_4_R0_en),
    .W0_addr(mem_113_4_W0_addr),
    .W0_clk(mem_113_4_W0_clk),
    .W0_data(mem_113_4_W0_data),
    .W0_en(mem_113_4_W0_en),
    .W0_mask(mem_113_4_W0_mask)
  );
  split_mem_0_ext mem_113_5 (
    .R0_addr(mem_113_5_R0_addr),
    .R0_clk(mem_113_5_R0_clk),
    .R0_data(mem_113_5_R0_data),
    .R0_en(mem_113_5_R0_en),
    .W0_addr(mem_113_5_W0_addr),
    .W0_clk(mem_113_5_W0_clk),
    .W0_data(mem_113_5_W0_data),
    .W0_en(mem_113_5_W0_en),
    .W0_mask(mem_113_5_W0_mask)
  );
  split_mem_0_ext mem_113_6 (
    .R0_addr(mem_113_6_R0_addr),
    .R0_clk(mem_113_6_R0_clk),
    .R0_data(mem_113_6_R0_data),
    .R0_en(mem_113_6_R0_en),
    .W0_addr(mem_113_6_W0_addr),
    .W0_clk(mem_113_6_W0_clk),
    .W0_data(mem_113_6_W0_data),
    .W0_en(mem_113_6_W0_en),
    .W0_mask(mem_113_6_W0_mask)
  );
  split_mem_0_ext mem_113_7 (
    .R0_addr(mem_113_7_R0_addr),
    .R0_clk(mem_113_7_R0_clk),
    .R0_data(mem_113_7_R0_data),
    .R0_en(mem_113_7_R0_en),
    .W0_addr(mem_113_7_W0_addr),
    .W0_clk(mem_113_7_W0_clk),
    .W0_data(mem_113_7_W0_data),
    .W0_en(mem_113_7_W0_en),
    .W0_mask(mem_113_7_W0_mask)
  );
  split_mem_0_ext mem_114_0 (
    .R0_addr(mem_114_0_R0_addr),
    .R0_clk(mem_114_0_R0_clk),
    .R0_data(mem_114_0_R0_data),
    .R0_en(mem_114_0_R0_en),
    .W0_addr(mem_114_0_W0_addr),
    .W0_clk(mem_114_0_W0_clk),
    .W0_data(mem_114_0_W0_data),
    .W0_en(mem_114_0_W0_en),
    .W0_mask(mem_114_0_W0_mask)
  );
  split_mem_0_ext mem_114_1 (
    .R0_addr(mem_114_1_R0_addr),
    .R0_clk(mem_114_1_R0_clk),
    .R0_data(mem_114_1_R0_data),
    .R0_en(mem_114_1_R0_en),
    .W0_addr(mem_114_1_W0_addr),
    .W0_clk(mem_114_1_W0_clk),
    .W0_data(mem_114_1_W0_data),
    .W0_en(mem_114_1_W0_en),
    .W0_mask(mem_114_1_W0_mask)
  );
  split_mem_0_ext mem_114_2 (
    .R0_addr(mem_114_2_R0_addr),
    .R0_clk(mem_114_2_R0_clk),
    .R0_data(mem_114_2_R0_data),
    .R0_en(mem_114_2_R0_en),
    .W0_addr(mem_114_2_W0_addr),
    .W0_clk(mem_114_2_W0_clk),
    .W0_data(mem_114_2_W0_data),
    .W0_en(mem_114_2_W0_en),
    .W0_mask(mem_114_2_W0_mask)
  );
  split_mem_0_ext mem_114_3 (
    .R0_addr(mem_114_3_R0_addr),
    .R0_clk(mem_114_3_R0_clk),
    .R0_data(mem_114_3_R0_data),
    .R0_en(mem_114_3_R0_en),
    .W0_addr(mem_114_3_W0_addr),
    .W0_clk(mem_114_3_W0_clk),
    .W0_data(mem_114_3_W0_data),
    .W0_en(mem_114_3_W0_en),
    .W0_mask(mem_114_3_W0_mask)
  );
  split_mem_0_ext mem_114_4 (
    .R0_addr(mem_114_4_R0_addr),
    .R0_clk(mem_114_4_R0_clk),
    .R0_data(mem_114_4_R0_data),
    .R0_en(mem_114_4_R0_en),
    .W0_addr(mem_114_4_W0_addr),
    .W0_clk(mem_114_4_W0_clk),
    .W0_data(mem_114_4_W0_data),
    .W0_en(mem_114_4_W0_en),
    .W0_mask(mem_114_4_W0_mask)
  );
  split_mem_0_ext mem_114_5 (
    .R0_addr(mem_114_5_R0_addr),
    .R0_clk(mem_114_5_R0_clk),
    .R0_data(mem_114_5_R0_data),
    .R0_en(mem_114_5_R0_en),
    .W0_addr(mem_114_5_W0_addr),
    .W0_clk(mem_114_5_W0_clk),
    .W0_data(mem_114_5_W0_data),
    .W0_en(mem_114_5_W0_en),
    .W0_mask(mem_114_5_W0_mask)
  );
  split_mem_0_ext mem_114_6 (
    .R0_addr(mem_114_6_R0_addr),
    .R0_clk(mem_114_6_R0_clk),
    .R0_data(mem_114_6_R0_data),
    .R0_en(mem_114_6_R0_en),
    .W0_addr(mem_114_6_W0_addr),
    .W0_clk(mem_114_6_W0_clk),
    .W0_data(mem_114_6_W0_data),
    .W0_en(mem_114_6_W0_en),
    .W0_mask(mem_114_6_W0_mask)
  );
  split_mem_0_ext mem_114_7 (
    .R0_addr(mem_114_7_R0_addr),
    .R0_clk(mem_114_7_R0_clk),
    .R0_data(mem_114_7_R0_data),
    .R0_en(mem_114_7_R0_en),
    .W0_addr(mem_114_7_W0_addr),
    .W0_clk(mem_114_7_W0_clk),
    .W0_data(mem_114_7_W0_data),
    .W0_en(mem_114_7_W0_en),
    .W0_mask(mem_114_7_W0_mask)
  );
  split_mem_0_ext mem_115_0 (
    .R0_addr(mem_115_0_R0_addr),
    .R0_clk(mem_115_0_R0_clk),
    .R0_data(mem_115_0_R0_data),
    .R0_en(mem_115_0_R0_en),
    .W0_addr(mem_115_0_W0_addr),
    .W0_clk(mem_115_0_W0_clk),
    .W0_data(mem_115_0_W0_data),
    .W0_en(mem_115_0_W0_en),
    .W0_mask(mem_115_0_W0_mask)
  );
  split_mem_0_ext mem_115_1 (
    .R0_addr(mem_115_1_R0_addr),
    .R0_clk(mem_115_1_R0_clk),
    .R0_data(mem_115_1_R0_data),
    .R0_en(mem_115_1_R0_en),
    .W0_addr(mem_115_1_W0_addr),
    .W0_clk(mem_115_1_W0_clk),
    .W0_data(mem_115_1_W0_data),
    .W0_en(mem_115_1_W0_en),
    .W0_mask(mem_115_1_W0_mask)
  );
  split_mem_0_ext mem_115_2 (
    .R0_addr(mem_115_2_R0_addr),
    .R0_clk(mem_115_2_R0_clk),
    .R0_data(mem_115_2_R0_data),
    .R0_en(mem_115_2_R0_en),
    .W0_addr(mem_115_2_W0_addr),
    .W0_clk(mem_115_2_W0_clk),
    .W0_data(mem_115_2_W0_data),
    .W0_en(mem_115_2_W0_en),
    .W0_mask(mem_115_2_W0_mask)
  );
  split_mem_0_ext mem_115_3 (
    .R0_addr(mem_115_3_R0_addr),
    .R0_clk(mem_115_3_R0_clk),
    .R0_data(mem_115_3_R0_data),
    .R0_en(mem_115_3_R0_en),
    .W0_addr(mem_115_3_W0_addr),
    .W0_clk(mem_115_3_W0_clk),
    .W0_data(mem_115_3_W0_data),
    .W0_en(mem_115_3_W0_en),
    .W0_mask(mem_115_3_W0_mask)
  );
  split_mem_0_ext mem_115_4 (
    .R0_addr(mem_115_4_R0_addr),
    .R0_clk(mem_115_4_R0_clk),
    .R0_data(mem_115_4_R0_data),
    .R0_en(mem_115_4_R0_en),
    .W0_addr(mem_115_4_W0_addr),
    .W0_clk(mem_115_4_W0_clk),
    .W0_data(mem_115_4_W0_data),
    .W0_en(mem_115_4_W0_en),
    .W0_mask(mem_115_4_W0_mask)
  );
  split_mem_0_ext mem_115_5 (
    .R0_addr(mem_115_5_R0_addr),
    .R0_clk(mem_115_5_R0_clk),
    .R0_data(mem_115_5_R0_data),
    .R0_en(mem_115_5_R0_en),
    .W0_addr(mem_115_5_W0_addr),
    .W0_clk(mem_115_5_W0_clk),
    .W0_data(mem_115_5_W0_data),
    .W0_en(mem_115_5_W0_en),
    .W0_mask(mem_115_5_W0_mask)
  );
  split_mem_0_ext mem_115_6 (
    .R0_addr(mem_115_6_R0_addr),
    .R0_clk(mem_115_6_R0_clk),
    .R0_data(mem_115_6_R0_data),
    .R0_en(mem_115_6_R0_en),
    .W0_addr(mem_115_6_W0_addr),
    .W0_clk(mem_115_6_W0_clk),
    .W0_data(mem_115_6_W0_data),
    .W0_en(mem_115_6_W0_en),
    .W0_mask(mem_115_6_W0_mask)
  );
  split_mem_0_ext mem_115_7 (
    .R0_addr(mem_115_7_R0_addr),
    .R0_clk(mem_115_7_R0_clk),
    .R0_data(mem_115_7_R0_data),
    .R0_en(mem_115_7_R0_en),
    .W0_addr(mem_115_7_W0_addr),
    .W0_clk(mem_115_7_W0_clk),
    .W0_data(mem_115_7_W0_data),
    .W0_en(mem_115_7_W0_en),
    .W0_mask(mem_115_7_W0_mask)
  );
  split_mem_0_ext mem_116_0 (
    .R0_addr(mem_116_0_R0_addr),
    .R0_clk(mem_116_0_R0_clk),
    .R0_data(mem_116_0_R0_data),
    .R0_en(mem_116_0_R0_en),
    .W0_addr(mem_116_0_W0_addr),
    .W0_clk(mem_116_0_W0_clk),
    .W0_data(mem_116_0_W0_data),
    .W0_en(mem_116_0_W0_en),
    .W0_mask(mem_116_0_W0_mask)
  );
  split_mem_0_ext mem_116_1 (
    .R0_addr(mem_116_1_R0_addr),
    .R0_clk(mem_116_1_R0_clk),
    .R0_data(mem_116_1_R0_data),
    .R0_en(mem_116_1_R0_en),
    .W0_addr(mem_116_1_W0_addr),
    .W0_clk(mem_116_1_W0_clk),
    .W0_data(mem_116_1_W0_data),
    .W0_en(mem_116_1_W0_en),
    .W0_mask(mem_116_1_W0_mask)
  );
  split_mem_0_ext mem_116_2 (
    .R0_addr(mem_116_2_R0_addr),
    .R0_clk(mem_116_2_R0_clk),
    .R0_data(mem_116_2_R0_data),
    .R0_en(mem_116_2_R0_en),
    .W0_addr(mem_116_2_W0_addr),
    .W0_clk(mem_116_2_W0_clk),
    .W0_data(mem_116_2_W0_data),
    .W0_en(mem_116_2_W0_en),
    .W0_mask(mem_116_2_W0_mask)
  );
  split_mem_0_ext mem_116_3 (
    .R0_addr(mem_116_3_R0_addr),
    .R0_clk(mem_116_3_R0_clk),
    .R0_data(mem_116_3_R0_data),
    .R0_en(mem_116_3_R0_en),
    .W0_addr(mem_116_3_W0_addr),
    .W0_clk(mem_116_3_W0_clk),
    .W0_data(mem_116_3_W0_data),
    .W0_en(mem_116_3_W0_en),
    .W0_mask(mem_116_3_W0_mask)
  );
  split_mem_0_ext mem_116_4 (
    .R0_addr(mem_116_4_R0_addr),
    .R0_clk(mem_116_4_R0_clk),
    .R0_data(mem_116_4_R0_data),
    .R0_en(mem_116_4_R0_en),
    .W0_addr(mem_116_4_W0_addr),
    .W0_clk(mem_116_4_W0_clk),
    .W0_data(mem_116_4_W0_data),
    .W0_en(mem_116_4_W0_en),
    .W0_mask(mem_116_4_W0_mask)
  );
  split_mem_0_ext mem_116_5 (
    .R0_addr(mem_116_5_R0_addr),
    .R0_clk(mem_116_5_R0_clk),
    .R0_data(mem_116_5_R0_data),
    .R0_en(mem_116_5_R0_en),
    .W0_addr(mem_116_5_W0_addr),
    .W0_clk(mem_116_5_W0_clk),
    .W0_data(mem_116_5_W0_data),
    .W0_en(mem_116_5_W0_en),
    .W0_mask(mem_116_5_W0_mask)
  );
  split_mem_0_ext mem_116_6 (
    .R0_addr(mem_116_6_R0_addr),
    .R0_clk(mem_116_6_R0_clk),
    .R0_data(mem_116_6_R0_data),
    .R0_en(mem_116_6_R0_en),
    .W0_addr(mem_116_6_W0_addr),
    .W0_clk(mem_116_6_W0_clk),
    .W0_data(mem_116_6_W0_data),
    .W0_en(mem_116_6_W0_en),
    .W0_mask(mem_116_6_W0_mask)
  );
  split_mem_0_ext mem_116_7 (
    .R0_addr(mem_116_7_R0_addr),
    .R0_clk(mem_116_7_R0_clk),
    .R0_data(mem_116_7_R0_data),
    .R0_en(mem_116_7_R0_en),
    .W0_addr(mem_116_7_W0_addr),
    .W0_clk(mem_116_7_W0_clk),
    .W0_data(mem_116_7_W0_data),
    .W0_en(mem_116_7_W0_en),
    .W0_mask(mem_116_7_W0_mask)
  );
  split_mem_0_ext mem_117_0 (
    .R0_addr(mem_117_0_R0_addr),
    .R0_clk(mem_117_0_R0_clk),
    .R0_data(mem_117_0_R0_data),
    .R0_en(mem_117_0_R0_en),
    .W0_addr(mem_117_0_W0_addr),
    .W0_clk(mem_117_0_W0_clk),
    .W0_data(mem_117_0_W0_data),
    .W0_en(mem_117_0_W0_en),
    .W0_mask(mem_117_0_W0_mask)
  );
  split_mem_0_ext mem_117_1 (
    .R0_addr(mem_117_1_R0_addr),
    .R0_clk(mem_117_1_R0_clk),
    .R0_data(mem_117_1_R0_data),
    .R0_en(mem_117_1_R0_en),
    .W0_addr(mem_117_1_W0_addr),
    .W0_clk(mem_117_1_W0_clk),
    .W0_data(mem_117_1_W0_data),
    .W0_en(mem_117_1_W0_en),
    .W0_mask(mem_117_1_W0_mask)
  );
  split_mem_0_ext mem_117_2 (
    .R0_addr(mem_117_2_R0_addr),
    .R0_clk(mem_117_2_R0_clk),
    .R0_data(mem_117_2_R0_data),
    .R0_en(mem_117_2_R0_en),
    .W0_addr(mem_117_2_W0_addr),
    .W0_clk(mem_117_2_W0_clk),
    .W0_data(mem_117_2_W0_data),
    .W0_en(mem_117_2_W0_en),
    .W0_mask(mem_117_2_W0_mask)
  );
  split_mem_0_ext mem_117_3 (
    .R0_addr(mem_117_3_R0_addr),
    .R0_clk(mem_117_3_R0_clk),
    .R0_data(mem_117_3_R0_data),
    .R0_en(mem_117_3_R0_en),
    .W0_addr(mem_117_3_W0_addr),
    .W0_clk(mem_117_3_W0_clk),
    .W0_data(mem_117_3_W0_data),
    .W0_en(mem_117_3_W0_en),
    .W0_mask(mem_117_3_W0_mask)
  );
  split_mem_0_ext mem_117_4 (
    .R0_addr(mem_117_4_R0_addr),
    .R0_clk(mem_117_4_R0_clk),
    .R0_data(mem_117_4_R0_data),
    .R0_en(mem_117_4_R0_en),
    .W0_addr(mem_117_4_W0_addr),
    .W0_clk(mem_117_4_W0_clk),
    .W0_data(mem_117_4_W0_data),
    .W0_en(mem_117_4_W0_en),
    .W0_mask(mem_117_4_W0_mask)
  );
  split_mem_0_ext mem_117_5 (
    .R0_addr(mem_117_5_R0_addr),
    .R0_clk(mem_117_5_R0_clk),
    .R0_data(mem_117_5_R0_data),
    .R0_en(mem_117_5_R0_en),
    .W0_addr(mem_117_5_W0_addr),
    .W0_clk(mem_117_5_W0_clk),
    .W0_data(mem_117_5_W0_data),
    .W0_en(mem_117_5_W0_en),
    .W0_mask(mem_117_5_W0_mask)
  );
  split_mem_0_ext mem_117_6 (
    .R0_addr(mem_117_6_R0_addr),
    .R0_clk(mem_117_6_R0_clk),
    .R0_data(mem_117_6_R0_data),
    .R0_en(mem_117_6_R0_en),
    .W0_addr(mem_117_6_W0_addr),
    .W0_clk(mem_117_6_W0_clk),
    .W0_data(mem_117_6_W0_data),
    .W0_en(mem_117_6_W0_en),
    .W0_mask(mem_117_6_W0_mask)
  );
  split_mem_0_ext mem_117_7 (
    .R0_addr(mem_117_7_R0_addr),
    .R0_clk(mem_117_7_R0_clk),
    .R0_data(mem_117_7_R0_data),
    .R0_en(mem_117_7_R0_en),
    .W0_addr(mem_117_7_W0_addr),
    .W0_clk(mem_117_7_W0_clk),
    .W0_data(mem_117_7_W0_data),
    .W0_en(mem_117_7_W0_en),
    .W0_mask(mem_117_7_W0_mask)
  );
  split_mem_0_ext mem_118_0 (
    .R0_addr(mem_118_0_R0_addr),
    .R0_clk(mem_118_0_R0_clk),
    .R0_data(mem_118_0_R0_data),
    .R0_en(mem_118_0_R0_en),
    .W0_addr(mem_118_0_W0_addr),
    .W0_clk(mem_118_0_W0_clk),
    .W0_data(mem_118_0_W0_data),
    .W0_en(mem_118_0_W0_en),
    .W0_mask(mem_118_0_W0_mask)
  );
  split_mem_0_ext mem_118_1 (
    .R0_addr(mem_118_1_R0_addr),
    .R0_clk(mem_118_1_R0_clk),
    .R0_data(mem_118_1_R0_data),
    .R0_en(mem_118_1_R0_en),
    .W0_addr(mem_118_1_W0_addr),
    .W0_clk(mem_118_1_W0_clk),
    .W0_data(mem_118_1_W0_data),
    .W0_en(mem_118_1_W0_en),
    .W0_mask(mem_118_1_W0_mask)
  );
  split_mem_0_ext mem_118_2 (
    .R0_addr(mem_118_2_R0_addr),
    .R0_clk(mem_118_2_R0_clk),
    .R0_data(mem_118_2_R0_data),
    .R0_en(mem_118_2_R0_en),
    .W0_addr(mem_118_2_W0_addr),
    .W0_clk(mem_118_2_W0_clk),
    .W0_data(mem_118_2_W0_data),
    .W0_en(mem_118_2_W0_en),
    .W0_mask(mem_118_2_W0_mask)
  );
  split_mem_0_ext mem_118_3 (
    .R0_addr(mem_118_3_R0_addr),
    .R0_clk(mem_118_3_R0_clk),
    .R0_data(mem_118_3_R0_data),
    .R0_en(mem_118_3_R0_en),
    .W0_addr(mem_118_3_W0_addr),
    .W0_clk(mem_118_3_W0_clk),
    .W0_data(mem_118_3_W0_data),
    .W0_en(mem_118_3_W0_en),
    .W0_mask(mem_118_3_W0_mask)
  );
  split_mem_0_ext mem_118_4 (
    .R0_addr(mem_118_4_R0_addr),
    .R0_clk(mem_118_4_R0_clk),
    .R0_data(mem_118_4_R0_data),
    .R0_en(mem_118_4_R0_en),
    .W0_addr(mem_118_4_W0_addr),
    .W0_clk(mem_118_4_W0_clk),
    .W0_data(mem_118_4_W0_data),
    .W0_en(mem_118_4_W0_en),
    .W0_mask(mem_118_4_W0_mask)
  );
  split_mem_0_ext mem_118_5 (
    .R0_addr(mem_118_5_R0_addr),
    .R0_clk(mem_118_5_R0_clk),
    .R0_data(mem_118_5_R0_data),
    .R0_en(mem_118_5_R0_en),
    .W0_addr(mem_118_5_W0_addr),
    .W0_clk(mem_118_5_W0_clk),
    .W0_data(mem_118_5_W0_data),
    .W0_en(mem_118_5_W0_en),
    .W0_mask(mem_118_5_W0_mask)
  );
  split_mem_0_ext mem_118_6 (
    .R0_addr(mem_118_6_R0_addr),
    .R0_clk(mem_118_6_R0_clk),
    .R0_data(mem_118_6_R0_data),
    .R0_en(mem_118_6_R0_en),
    .W0_addr(mem_118_6_W0_addr),
    .W0_clk(mem_118_6_W0_clk),
    .W0_data(mem_118_6_W0_data),
    .W0_en(mem_118_6_W0_en),
    .W0_mask(mem_118_6_W0_mask)
  );
  split_mem_0_ext mem_118_7 (
    .R0_addr(mem_118_7_R0_addr),
    .R0_clk(mem_118_7_R0_clk),
    .R0_data(mem_118_7_R0_data),
    .R0_en(mem_118_7_R0_en),
    .W0_addr(mem_118_7_W0_addr),
    .W0_clk(mem_118_7_W0_clk),
    .W0_data(mem_118_7_W0_data),
    .W0_en(mem_118_7_W0_en),
    .W0_mask(mem_118_7_W0_mask)
  );
  split_mem_0_ext mem_119_0 (
    .R0_addr(mem_119_0_R0_addr),
    .R0_clk(mem_119_0_R0_clk),
    .R0_data(mem_119_0_R0_data),
    .R0_en(mem_119_0_R0_en),
    .W0_addr(mem_119_0_W0_addr),
    .W0_clk(mem_119_0_W0_clk),
    .W0_data(mem_119_0_W0_data),
    .W0_en(mem_119_0_W0_en),
    .W0_mask(mem_119_0_W0_mask)
  );
  split_mem_0_ext mem_119_1 (
    .R0_addr(mem_119_1_R0_addr),
    .R0_clk(mem_119_1_R0_clk),
    .R0_data(mem_119_1_R0_data),
    .R0_en(mem_119_1_R0_en),
    .W0_addr(mem_119_1_W0_addr),
    .W0_clk(mem_119_1_W0_clk),
    .W0_data(mem_119_1_W0_data),
    .W0_en(mem_119_1_W0_en),
    .W0_mask(mem_119_1_W0_mask)
  );
  split_mem_0_ext mem_119_2 (
    .R0_addr(mem_119_2_R0_addr),
    .R0_clk(mem_119_2_R0_clk),
    .R0_data(mem_119_2_R0_data),
    .R0_en(mem_119_2_R0_en),
    .W0_addr(mem_119_2_W0_addr),
    .W0_clk(mem_119_2_W0_clk),
    .W0_data(mem_119_2_W0_data),
    .W0_en(mem_119_2_W0_en),
    .W0_mask(mem_119_2_W0_mask)
  );
  split_mem_0_ext mem_119_3 (
    .R0_addr(mem_119_3_R0_addr),
    .R0_clk(mem_119_3_R0_clk),
    .R0_data(mem_119_3_R0_data),
    .R0_en(mem_119_3_R0_en),
    .W0_addr(mem_119_3_W0_addr),
    .W0_clk(mem_119_3_W0_clk),
    .W0_data(mem_119_3_W0_data),
    .W0_en(mem_119_3_W0_en),
    .W0_mask(mem_119_3_W0_mask)
  );
  split_mem_0_ext mem_119_4 (
    .R0_addr(mem_119_4_R0_addr),
    .R0_clk(mem_119_4_R0_clk),
    .R0_data(mem_119_4_R0_data),
    .R0_en(mem_119_4_R0_en),
    .W0_addr(mem_119_4_W0_addr),
    .W0_clk(mem_119_4_W0_clk),
    .W0_data(mem_119_4_W0_data),
    .W0_en(mem_119_4_W0_en),
    .W0_mask(mem_119_4_W0_mask)
  );
  split_mem_0_ext mem_119_5 (
    .R0_addr(mem_119_5_R0_addr),
    .R0_clk(mem_119_5_R0_clk),
    .R0_data(mem_119_5_R0_data),
    .R0_en(mem_119_5_R0_en),
    .W0_addr(mem_119_5_W0_addr),
    .W0_clk(mem_119_5_W0_clk),
    .W0_data(mem_119_5_W0_data),
    .W0_en(mem_119_5_W0_en),
    .W0_mask(mem_119_5_W0_mask)
  );
  split_mem_0_ext mem_119_6 (
    .R0_addr(mem_119_6_R0_addr),
    .R0_clk(mem_119_6_R0_clk),
    .R0_data(mem_119_6_R0_data),
    .R0_en(mem_119_6_R0_en),
    .W0_addr(mem_119_6_W0_addr),
    .W0_clk(mem_119_6_W0_clk),
    .W0_data(mem_119_6_W0_data),
    .W0_en(mem_119_6_W0_en),
    .W0_mask(mem_119_6_W0_mask)
  );
  split_mem_0_ext mem_119_7 (
    .R0_addr(mem_119_7_R0_addr),
    .R0_clk(mem_119_7_R0_clk),
    .R0_data(mem_119_7_R0_data),
    .R0_en(mem_119_7_R0_en),
    .W0_addr(mem_119_7_W0_addr),
    .W0_clk(mem_119_7_W0_clk),
    .W0_data(mem_119_7_W0_data),
    .W0_en(mem_119_7_W0_en),
    .W0_mask(mem_119_7_W0_mask)
  );
  split_mem_0_ext mem_120_0 (
    .R0_addr(mem_120_0_R0_addr),
    .R0_clk(mem_120_0_R0_clk),
    .R0_data(mem_120_0_R0_data),
    .R0_en(mem_120_0_R0_en),
    .W0_addr(mem_120_0_W0_addr),
    .W0_clk(mem_120_0_W0_clk),
    .W0_data(mem_120_0_W0_data),
    .W0_en(mem_120_0_W0_en),
    .W0_mask(mem_120_0_W0_mask)
  );
  split_mem_0_ext mem_120_1 (
    .R0_addr(mem_120_1_R0_addr),
    .R0_clk(mem_120_1_R0_clk),
    .R0_data(mem_120_1_R0_data),
    .R0_en(mem_120_1_R0_en),
    .W0_addr(mem_120_1_W0_addr),
    .W0_clk(mem_120_1_W0_clk),
    .W0_data(mem_120_1_W0_data),
    .W0_en(mem_120_1_W0_en),
    .W0_mask(mem_120_1_W0_mask)
  );
  split_mem_0_ext mem_120_2 (
    .R0_addr(mem_120_2_R0_addr),
    .R0_clk(mem_120_2_R0_clk),
    .R0_data(mem_120_2_R0_data),
    .R0_en(mem_120_2_R0_en),
    .W0_addr(mem_120_2_W0_addr),
    .W0_clk(mem_120_2_W0_clk),
    .W0_data(mem_120_2_W0_data),
    .W0_en(mem_120_2_W0_en),
    .W0_mask(mem_120_2_W0_mask)
  );
  split_mem_0_ext mem_120_3 (
    .R0_addr(mem_120_3_R0_addr),
    .R0_clk(mem_120_3_R0_clk),
    .R0_data(mem_120_3_R0_data),
    .R0_en(mem_120_3_R0_en),
    .W0_addr(mem_120_3_W0_addr),
    .W0_clk(mem_120_3_W0_clk),
    .W0_data(mem_120_3_W0_data),
    .W0_en(mem_120_3_W0_en),
    .W0_mask(mem_120_3_W0_mask)
  );
  split_mem_0_ext mem_120_4 (
    .R0_addr(mem_120_4_R0_addr),
    .R0_clk(mem_120_4_R0_clk),
    .R0_data(mem_120_4_R0_data),
    .R0_en(mem_120_4_R0_en),
    .W0_addr(mem_120_4_W0_addr),
    .W0_clk(mem_120_4_W0_clk),
    .W0_data(mem_120_4_W0_data),
    .W0_en(mem_120_4_W0_en),
    .W0_mask(mem_120_4_W0_mask)
  );
  split_mem_0_ext mem_120_5 (
    .R0_addr(mem_120_5_R0_addr),
    .R0_clk(mem_120_5_R0_clk),
    .R0_data(mem_120_5_R0_data),
    .R0_en(mem_120_5_R0_en),
    .W0_addr(mem_120_5_W0_addr),
    .W0_clk(mem_120_5_W0_clk),
    .W0_data(mem_120_5_W0_data),
    .W0_en(mem_120_5_W0_en),
    .W0_mask(mem_120_5_W0_mask)
  );
  split_mem_0_ext mem_120_6 (
    .R0_addr(mem_120_6_R0_addr),
    .R0_clk(mem_120_6_R0_clk),
    .R0_data(mem_120_6_R0_data),
    .R0_en(mem_120_6_R0_en),
    .W0_addr(mem_120_6_W0_addr),
    .W0_clk(mem_120_6_W0_clk),
    .W0_data(mem_120_6_W0_data),
    .W0_en(mem_120_6_W0_en),
    .W0_mask(mem_120_6_W0_mask)
  );
  split_mem_0_ext mem_120_7 (
    .R0_addr(mem_120_7_R0_addr),
    .R0_clk(mem_120_7_R0_clk),
    .R0_data(mem_120_7_R0_data),
    .R0_en(mem_120_7_R0_en),
    .W0_addr(mem_120_7_W0_addr),
    .W0_clk(mem_120_7_W0_clk),
    .W0_data(mem_120_7_W0_data),
    .W0_en(mem_120_7_W0_en),
    .W0_mask(mem_120_7_W0_mask)
  );
  split_mem_0_ext mem_121_0 (
    .R0_addr(mem_121_0_R0_addr),
    .R0_clk(mem_121_0_R0_clk),
    .R0_data(mem_121_0_R0_data),
    .R0_en(mem_121_0_R0_en),
    .W0_addr(mem_121_0_W0_addr),
    .W0_clk(mem_121_0_W0_clk),
    .W0_data(mem_121_0_W0_data),
    .W0_en(mem_121_0_W0_en),
    .W0_mask(mem_121_0_W0_mask)
  );
  split_mem_0_ext mem_121_1 (
    .R0_addr(mem_121_1_R0_addr),
    .R0_clk(mem_121_1_R0_clk),
    .R0_data(mem_121_1_R0_data),
    .R0_en(mem_121_1_R0_en),
    .W0_addr(mem_121_1_W0_addr),
    .W0_clk(mem_121_1_W0_clk),
    .W0_data(mem_121_1_W0_data),
    .W0_en(mem_121_1_W0_en),
    .W0_mask(mem_121_1_W0_mask)
  );
  split_mem_0_ext mem_121_2 (
    .R0_addr(mem_121_2_R0_addr),
    .R0_clk(mem_121_2_R0_clk),
    .R0_data(mem_121_2_R0_data),
    .R0_en(mem_121_2_R0_en),
    .W0_addr(mem_121_2_W0_addr),
    .W0_clk(mem_121_2_W0_clk),
    .W0_data(mem_121_2_W0_data),
    .W0_en(mem_121_2_W0_en),
    .W0_mask(mem_121_2_W0_mask)
  );
  split_mem_0_ext mem_121_3 (
    .R0_addr(mem_121_3_R0_addr),
    .R0_clk(mem_121_3_R0_clk),
    .R0_data(mem_121_3_R0_data),
    .R0_en(mem_121_3_R0_en),
    .W0_addr(mem_121_3_W0_addr),
    .W0_clk(mem_121_3_W0_clk),
    .W0_data(mem_121_3_W0_data),
    .W0_en(mem_121_3_W0_en),
    .W0_mask(mem_121_3_W0_mask)
  );
  split_mem_0_ext mem_121_4 (
    .R0_addr(mem_121_4_R0_addr),
    .R0_clk(mem_121_4_R0_clk),
    .R0_data(mem_121_4_R0_data),
    .R0_en(mem_121_4_R0_en),
    .W0_addr(mem_121_4_W0_addr),
    .W0_clk(mem_121_4_W0_clk),
    .W0_data(mem_121_4_W0_data),
    .W0_en(mem_121_4_W0_en),
    .W0_mask(mem_121_4_W0_mask)
  );
  split_mem_0_ext mem_121_5 (
    .R0_addr(mem_121_5_R0_addr),
    .R0_clk(mem_121_5_R0_clk),
    .R0_data(mem_121_5_R0_data),
    .R0_en(mem_121_5_R0_en),
    .W0_addr(mem_121_5_W0_addr),
    .W0_clk(mem_121_5_W0_clk),
    .W0_data(mem_121_5_W0_data),
    .W0_en(mem_121_5_W0_en),
    .W0_mask(mem_121_5_W0_mask)
  );
  split_mem_0_ext mem_121_6 (
    .R0_addr(mem_121_6_R0_addr),
    .R0_clk(mem_121_6_R0_clk),
    .R0_data(mem_121_6_R0_data),
    .R0_en(mem_121_6_R0_en),
    .W0_addr(mem_121_6_W0_addr),
    .W0_clk(mem_121_6_W0_clk),
    .W0_data(mem_121_6_W0_data),
    .W0_en(mem_121_6_W0_en),
    .W0_mask(mem_121_6_W0_mask)
  );
  split_mem_0_ext mem_121_7 (
    .R0_addr(mem_121_7_R0_addr),
    .R0_clk(mem_121_7_R0_clk),
    .R0_data(mem_121_7_R0_data),
    .R0_en(mem_121_7_R0_en),
    .W0_addr(mem_121_7_W0_addr),
    .W0_clk(mem_121_7_W0_clk),
    .W0_data(mem_121_7_W0_data),
    .W0_en(mem_121_7_W0_en),
    .W0_mask(mem_121_7_W0_mask)
  );
  split_mem_0_ext mem_122_0 (
    .R0_addr(mem_122_0_R0_addr),
    .R0_clk(mem_122_0_R0_clk),
    .R0_data(mem_122_0_R0_data),
    .R0_en(mem_122_0_R0_en),
    .W0_addr(mem_122_0_W0_addr),
    .W0_clk(mem_122_0_W0_clk),
    .W0_data(mem_122_0_W0_data),
    .W0_en(mem_122_0_W0_en),
    .W0_mask(mem_122_0_W0_mask)
  );
  split_mem_0_ext mem_122_1 (
    .R0_addr(mem_122_1_R0_addr),
    .R0_clk(mem_122_1_R0_clk),
    .R0_data(mem_122_1_R0_data),
    .R0_en(mem_122_1_R0_en),
    .W0_addr(mem_122_1_W0_addr),
    .W0_clk(mem_122_1_W0_clk),
    .W0_data(mem_122_1_W0_data),
    .W0_en(mem_122_1_W0_en),
    .W0_mask(mem_122_1_W0_mask)
  );
  split_mem_0_ext mem_122_2 (
    .R0_addr(mem_122_2_R0_addr),
    .R0_clk(mem_122_2_R0_clk),
    .R0_data(mem_122_2_R0_data),
    .R0_en(mem_122_2_R0_en),
    .W0_addr(mem_122_2_W0_addr),
    .W0_clk(mem_122_2_W0_clk),
    .W0_data(mem_122_2_W0_data),
    .W0_en(mem_122_2_W0_en),
    .W0_mask(mem_122_2_W0_mask)
  );
  split_mem_0_ext mem_122_3 (
    .R0_addr(mem_122_3_R0_addr),
    .R0_clk(mem_122_3_R0_clk),
    .R0_data(mem_122_3_R0_data),
    .R0_en(mem_122_3_R0_en),
    .W0_addr(mem_122_3_W0_addr),
    .W0_clk(mem_122_3_W0_clk),
    .W0_data(mem_122_3_W0_data),
    .W0_en(mem_122_3_W0_en),
    .W0_mask(mem_122_3_W0_mask)
  );
  split_mem_0_ext mem_122_4 (
    .R0_addr(mem_122_4_R0_addr),
    .R0_clk(mem_122_4_R0_clk),
    .R0_data(mem_122_4_R0_data),
    .R0_en(mem_122_4_R0_en),
    .W0_addr(mem_122_4_W0_addr),
    .W0_clk(mem_122_4_W0_clk),
    .W0_data(mem_122_4_W0_data),
    .W0_en(mem_122_4_W0_en),
    .W0_mask(mem_122_4_W0_mask)
  );
  split_mem_0_ext mem_122_5 (
    .R0_addr(mem_122_5_R0_addr),
    .R0_clk(mem_122_5_R0_clk),
    .R0_data(mem_122_5_R0_data),
    .R0_en(mem_122_5_R0_en),
    .W0_addr(mem_122_5_W0_addr),
    .W0_clk(mem_122_5_W0_clk),
    .W0_data(mem_122_5_W0_data),
    .W0_en(mem_122_5_W0_en),
    .W0_mask(mem_122_5_W0_mask)
  );
  split_mem_0_ext mem_122_6 (
    .R0_addr(mem_122_6_R0_addr),
    .R0_clk(mem_122_6_R0_clk),
    .R0_data(mem_122_6_R0_data),
    .R0_en(mem_122_6_R0_en),
    .W0_addr(mem_122_6_W0_addr),
    .W0_clk(mem_122_6_W0_clk),
    .W0_data(mem_122_6_W0_data),
    .W0_en(mem_122_6_W0_en),
    .W0_mask(mem_122_6_W0_mask)
  );
  split_mem_0_ext mem_122_7 (
    .R0_addr(mem_122_7_R0_addr),
    .R0_clk(mem_122_7_R0_clk),
    .R0_data(mem_122_7_R0_data),
    .R0_en(mem_122_7_R0_en),
    .W0_addr(mem_122_7_W0_addr),
    .W0_clk(mem_122_7_W0_clk),
    .W0_data(mem_122_7_W0_data),
    .W0_en(mem_122_7_W0_en),
    .W0_mask(mem_122_7_W0_mask)
  );
  split_mem_0_ext mem_123_0 (
    .R0_addr(mem_123_0_R0_addr),
    .R0_clk(mem_123_0_R0_clk),
    .R0_data(mem_123_0_R0_data),
    .R0_en(mem_123_0_R0_en),
    .W0_addr(mem_123_0_W0_addr),
    .W0_clk(mem_123_0_W0_clk),
    .W0_data(mem_123_0_W0_data),
    .W0_en(mem_123_0_W0_en),
    .W0_mask(mem_123_0_W0_mask)
  );
  split_mem_0_ext mem_123_1 (
    .R0_addr(mem_123_1_R0_addr),
    .R0_clk(mem_123_1_R0_clk),
    .R0_data(mem_123_1_R0_data),
    .R0_en(mem_123_1_R0_en),
    .W0_addr(mem_123_1_W0_addr),
    .W0_clk(mem_123_1_W0_clk),
    .W0_data(mem_123_1_W0_data),
    .W0_en(mem_123_1_W0_en),
    .W0_mask(mem_123_1_W0_mask)
  );
  split_mem_0_ext mem_123_2 (
    .R0_addr(mem_123_2_R0_addr),
    .R0_clk(mem_123_2_R0_clk),
    .R0_data(mem_123_2_R0_data),
    .R0_en(mem_123_2_R0_en),
    .W0_addr(mem_123_2_W0_addr),
    .W0_clk(mem_123_2_W0_clk),
    .W0_data(mem_123_2_W0_data),
    .W0_en(mem_123_2_W0_en),
    .W0_mask(mem_123_2_W0_mask)
  );
  split_mem_0_ext mem_123_3 (
    .R0_addr(mem_123_3_R0_addr),
    .R0_clk(mem_123_3_R0_clk),
    .R0_data(mem_123_3_R0_data),
    .R0_en(mem_123_3_R0_en),
    .W0_addr(mem_123_3_W0_addr),
    .W0_clk(mem_123_3_W0_clk),
    .W0_data(mem_123_3_W0_data),
    .W0_en(mem_123_3_W0_en),
    .W0_mask(mem_123_3_W0_mask)
  );
  split_mem_0_ext mem_123_4 (
    .R0_addr(mem_123_4_R0_addr),
    .R0_clk(mem_123_4_R0_clk),
    .R0_data(mem_123_4_R0_data),
    .R0_en(mem_123_4_R0_en),
    .W0_addr(mem_123_4_W0_addr),
    .W0_clk(mem_123_4_W0_clk),
    .W0_data(mem_123_4_W0_data),
    .W0_en(mem_123_4_W0_en),
    .W0_mask(mem_123_4_W0_mask)
  );
  split_mem_0_ext mem_123_5 (
    .R0_addr(mem_123_5_R0_addr),
    .R0_clk(mem_123_5_R0_clk),
    .R0_data(mem_123_5_R0_data),
    .R0_en(mem_123_5_R0_en),
    .W0_addr(mem_123_5_W0_addr),
    .W0_clk(mem_123_5_W0_clk),
    .W0_data(mem_123_5_W0_data),
    .W0_en(mem_123_5_W0_en),
    .W0_mask(mem_123_5_W0_mask)
  );
  split_mem_0_ext mem_123_6 (
    .R0_addr(mem_123_6_R0_addr),
    .R0_clk(mem_123_6_R0_clk),
    .R0_data(mem_123_6_R0_data),
    .R0_en(mem_123_6_R0_en),
    .W0_addr(mem_123_6_W0_addr),
    .W0_clk(mem_123_6_W0_clk),
    .W0_data(mem_123_6_W0_data),
    .W0_en(mem_123_6_W0_en),
    .W0_mask(mem_123_6_W0_mask)
  );
  split_mem_0_ext mem_123_7 (
    .R0_addr(mem_123_7_R0_addr),
    .R0_clk(mem_123_7_R0_clk),
    .R0_data(mem_123_7_R0_data),
    .R0_en(mem_123_7_R0_en),
    .W0_addr(mem_123_7_W0_addr),
    .W0_clk(mem_123_7_W0_clk),
    .W0_data(mem_123_7_W0_data),
    .W0_en(mem_123_7_W0_en),
    .W0_mask(mem_123_7_W0_mask)
  );
  split_mem_0_ext mem_124_0 (
    .R0_addr(mem_124_0_R0_addr),
    .R0_clk(mem_124_0_R0_clk),
    .R0_data(mem_124_0_R0_data),
    .R0_en(mem_124_0_R0_en),
    .W0_addr(mem_124_0_W0_addr),
    .W0_clk(mem_124_0_W0_clk),
    .W0_data(mem_124_0_W0_data),
    .W0_en(mem_124_0_W0_en),
    .W0_mask(mem_124_0_W0_mask)
  );
  split_mem_0_ext mem_124_1 (
    .R0_addr(mem_124_1_R0_addr),
    .R0_clk(mem_124_1_R0_clk),
    .R0_data(mem_124_1_R0_data),
    .R0_en(mem_124_1_R0_en),
    .W0_addr(mem_124_1_W0_addr),
    .W0_clk(mem_124_1_W0_clk),
    .W0_data(mem_124_1_W0_data),
    .W0_en(mem_124_1_W0_en),
    .W0_mask(mem_124_1_W0_mask)
  );
  split_mem_0_ext mem_124_2 (
    .R0_addr(mem_124_2_R0_addr),
    .R0_clk(mem_124_2_R0_clk),
    .R0_data(mem_124_2_R0_data),
    .R0_en(mem_124_2_R0_en),
    .W0_addr(mem_124_2_W0_addr),
    .W0_clk(mem_124_2_W0_clk),
    .W0_data(mem_124_2_W0_data),
    .W0_en(mem_124_2_W0_en),
    .W0_mask(mem_124_2_W0_mask)
  );
  split_mem_0_ext mem_124_3 (
    .R0_addr(mem_124_3_R0_addr),
    .R0_clk(mem_124_3_R0_clk),
    .R0_data(mem_124_3_R0_data),
    .R0_en(mem_124_3_R0_en),
    .W0_addr(mem_124_3_W0_addr),
    .W0_clk(mem_124_3_W0_clk),
    .W0_data(mem_124_3_W0_data),
    .W0_en(mem_124_3_W0_en),
    .W0_mask(mem_124_3_W0_mask)
  );
  split_mem_0_ext mem_124_4 (
    .R0_addr(mem_124_4_R0_addr),
    .R0_clk(mem_124_4_R0_clk),
    .R0_data(mem_124_4_R0_data),
    .R0_en(mem_124_4_R0_en),
    .W0_addr(mem_124_4_W0_addr),
    .W0_clk(mem_124_4_W0_clk),
    .W0_data(mem_124_4_W0_data),
    .W0_en(mem_124_4_W0_en),
    .W0_mask(mem_124_4_W0_mask)
  );
  split_mem_0_ext mem_124_5 (
    .R0_addr(mem_124_5_R0_addr),
    .R0_clk(mem_124_5_R0_clk),
    .R0_data(mem_124_5_R0_data),
    .R0_en(mem_124_5_R0_en),
    .W0_addr(mem_124_5_W0_addr),
    .W0_clk(mem_124_5_W0_clk),
    .W0_data(mem_124_5_W0_data),
    .W0_en(mem_124_5_W0_en),
    .W0_mask(mem_124_5_W0_mask)
  );
  split_mem_0_ext mem_124_6 (
    .R0_addr(mem_124_6_R0_addr),
    .R0_clk(mem_124_6_R0_clk),
    .R0_data(mem_124_6_R0_data),
    .R0_en(mem_124_6_R0_en),
    .W0_addr(mem_124_6_W0_addr),
    .W0_clk(mem_124_6_W0_clk),
    .W0_data(mem_124_6_W0_data),
    .W0_en(mem_124_6_W0_en),
    .W0_mask(mem_124_6_W0_mask)
  );
  split_mem_0_ext mem_124_7 (
    .R0_addr(mem_124_7_R0_addr),
    .R0_clk(mem_124_7_R0_clk),
    .R0_data(mem_124_7_R0_data),
    .R0_en(mem_124_7_R0_en),
    .W0_addr(mem_124_7_W0_addr),
    .W0_clk(mem_124_7_W0_clk),
    .W0_data(mem_124_7_W0_data),
    .W0_en(mem_124_7_W0_en),
    .W0_mask(mem_124_7_W0_mask)
  );
  split_mem_0_ext mem_125_0 (
    .R0_addr(mem_125_0_R0_addr),
    .R0_clk(mem_125_0_R0_clk),
    .R0_data(mem_125_0_R0_data),
    .R0_en(mem_125_0_R0_en),
    .W0_addr(mem_125_0_W0_addr),
    .W0_clk(mem_125_0_W0_clk),
    .W0_data(mem_125_0_W0_data),
    .W0_en(mem_125_0_W0_en),
    .W0_mask(mem_125_0_W0_mask)
  );
  split_mem_0_ext mem_125_1 (
    .R0_addr(mem_125_1_R0_addr),
    .R0_clk(mem_125_1_R0_clk),
    .R0_data(mem_125_1_R0_data),
    .R0_en(mem_125_1_R0_en),
    .W0_addr(mem_125_1_W0_addr),
    .W0_clk(mem_125_1_W0_clk),
    .W0_data(mem_125_1_W0_data),
    .W0_en(mem_125_1_W0_en),
    .W0_mask(mem_125_1_W0_mask)
  );
  split_mem_0_ext mem_125_2 (
    .R0_addr(mem_125_2_R0_addr),
    .R0_clk(mem_125_2_R0_clk),
    .R0_data(mem_125_2_R0_data),
    .R0_en(mem_125_2_R0_en),
    .W0_addr(mem_125_2_W0_addr),
    .W0_clk(mem_125_2_W0_clk),
    .W0_data(mem_125_2_W0_data),
    .W0_en(mem_125_2_W0_en),
    .W0_mask(mem_125_2_W0_mask)
  );
  split_mem_0_ext mem_125_3 (
    .R0_addr(mem_125_3_R0_addr),
    .R0_clk(mem_125_3_R0_clk),
    .R0_data(mem_125_3_R0_data),
    .R0_en(mem_125_3_R0_en),
    .W0_addr(mem_125_3_W0_addr),
    .W0_clk(mem_125_3_W0_clk),
    .W0_data(mem_125_3_W0_data),
    .W0_en(mem_125_3_W0_en),
    .W0_mask(mem_125_3_W0_mask)
  );
  split_mem_0_ext mem_125_4 (
    .R0_addr(mem_125_4_R0_addr),
    .R0_clk(mem_125_4_R0_clk),
    .R0_data(mem_125_4_R0_data),
    .R0_en(mem_125_4_R0_en),
    .W0_addr(mem_125_4_W0_addr),
    .W0_clk(mem_125_4_W0_clk),
    .W0_data(mem_125_4_W0_data),
    .W0_en(mem_125_4_W0_en),
    .W0_mask(mem_125_4_W0_mask)
  );
  split_mem_0_ext mem_125_5 (
    .R0_addr(mem_125_5_R0_addr),
    .R0_clk(mem_125_5_R0_clk),
    .R0_data(mem_125_5_R0_data),
    .R0_en(mem_125_5_R0_en),
    .W0_addr(mem_125_5_W0_addr),
    .W0_clk(mem_125_5_W0_clk),
    .W0_data(mem_125_5_W0_data),
    .W0_en(mem_125_5_W0_en),
    .W0_mask(mem_125_5_W0_mask)
  );
  split_mem_0_ext mem_125_6 (
    .R0_addr(mem_125_6_R0_addr),
    .R0_clk(mem_125_6_R0_clk),
    .R0_data(mem_125_6_R0_data),
    .R0_en(mem_125_6_R0_en),
    .W0_addr(mem_125_6_W0_addr),
    .W0_clk(mem_125_6_W0_clk),
    .W0_data(mem_125_6_W0_data),
    .W0_en(mem_125_6_W0_en),
    .W0_mask(mem_125_6_W0_mask)
  );
  split_mem_0_ext mem_125_7 (
    .R0_addr(mem_125_7_R0_addr),
    .R0_clk(mem_125_7_R0_clk),
    .R0_data(mem_125_7_R0_data),
    .R0_en(mem_125_7_R0_en),
    .W0_addr(mem_125_7_W0_addr),
    .W0_clk(mem_125_7_W0_clk),
    .W0_data(mem_125_7_W0_data),
    .W0_en(mem_125_7_W0_en),
    .W0_mask(mem_125_7_W0_mask)
  );
  split_mem_0_ext mem_126_0 (
    .R0_addr(mem_126_0_R0_addr),
    .R0_clk(mem_126_0_R0_clk),
    .R0_data(mem_126_0_R0_data),
    .R0_en(mem_126_0_R0_en),
    .W0_addr(mem_126_0_W0_addr),
    .W0_clk(mem_126_0_W0_clk),
    .W0_data(mem_126_0_W0_data),
    .W0_en(mem_126_0_W0_en),
    .W0_mask(mem_126_0_W0_mask)
  );
  split_mem_0_ext mem_126_1 (
    .R0_addr(mem_126_1_R0_addr),
    .R0_clk(mem_126_1_R0_clk),
    .R0_data(mem_126_1_R0_data),
    .R0_en(mem_126_1_R0_en),
    .W0_addr(mem_126_1_W0_addr),
    .W0_clk(mem_126_1_W0_clk),
    .W0_data(mem_126_1_W0_data),
    .W0_en(mem_126_1_W0_en),
    .W0_mask(mem_126_1_W0_mask)
  );
  split_mem_0_ext mem_126_2 (
    .R0_addr(mem_126_2_R0_addr),
    .R0_clk(mem_126_2_R0_clk),
    .R0_data(mem_126_2_R0_data),
    .R0_en(mem_126_2_R0_en),
    .W0_addr(mem_126_2_W0_addr),
    .W0_clk(mem_126_2_W0_clk),
    .W0_data(mem_126_2_W0_data),
    .W0_en(mem_126_2_W0_en),
    .W0_mask(mem_126_2_W0_mask)
  );
  split_mem_0_ext mem_126_3 (
    .R0_addr(mem_126_3_R0_addr),
    .R0_clk(mem_126_3_R0_clk),
    .R0_data(mem_126_3_R0_data),
    .R0_en(mem_126_3_R0_en),
    .W0_addr(mem_126_3_W0_addr),
    .W0_clk(mem_126_3_W0_clk),
    .W0_data(mem_126_3_W0_data),
    .W0_en(mem_126_3_W0_en),
    .W0_mask(mem_126_3_W0_mask)
  );
  split_mem_0_ext mem_126_4 (
    .R0_addr(mem_126_4_R0_addr),
    .R0_clk(mem_126_4_R0_clk),
    .R0_data(mem_126_4_R0_data),
    .R0_en(mem_126_4_R0_en),
    .W0_addr(mem_126_4_W0_addr),
    .W0_clk(mem_126_4_W0_clk),
    .W0_data(mem_126_4_W0_data),
    .W0_en(mem_126_4_W0_en),
    .W0_mask(mem_126_4_W0_mask)
  );
  split_mem_0_ext mem_126_5 (
    .R0_addr(mem_126_5_R0_addr),
    .R0_clk(mem_126_5_R0_clk),
    .R0_data(mem_126_5_R0_data),
    .R0_en(mem_126_5_R0_en),
    .W0_addr(mem_126_5_W0_addr),
    .W0_clk(mem_126_5_W0_clk),
    .W0_data(mem_126_5_W0_data),
    .W0_en(mem_126_5_W0_en),
    .W0_mask(mem_126_5_W0_mask)
  );
  split_mem_0_ext mem_126_6 (
    .R0_addr(mem_126_6_R0_addr),
    .R0_clk(mem_126_6_R0_clk),
    .R0_data(mem_126_6_R0_data),
    .R0_en(mem_126_6_R0_en),
    .W0_addr(mem_126_6_W0_addr),
    .W0_clk(mem_126_6_W0_clk),
    .W0_data(mem_126_6_W0_data),
    .W0_en(mem_126_6_W0_en),
    .W0_mask(mem_126_6_W0_mask)
  );
  split_mem_0_ext mem_126_7 (
    .R0_addr(mem_126_7_R0_addr),
    .R0_clk(mem_126_7_R0_clk),
    .R0_data(mem_126_7_R0_data),
    .R0_en(mem_126_7_R0_en),
    .W0_addr(mem_126_7_W0_addr),
    .W0_clk(mem_126_7_W0_clk),
    .W0_data(mem_126_7_W0_data),
    .W0_en(mem_126_7_W0_en),
    .W0_mask(mem_126_7_W0_mask)
  );
  split_mem_0_ext mem_127_0 (
    .R0_addr(mem_127_0_R0_addr),
    .R0_clk(mem_127_0_R0_clk),
    .R0_data(mem_127_0_R0_data),
    .R0_en(mem_127_0_R0_en),
    .W0_addr(mem_127_0_W0_addr),
    .W0_clk(mem_127_0_W0_clk),
    .W0_data(mem_127_0_W0_data),
    .W0_en(mem_127_0_W0_en),
    .W0_mask(mem_127_0_W0_mask)
  );
  split_mem_0_ext mem_127_1 (
    .R0_addr(mem_127_1_R0_addr),
    .R0_clk(mem_127_1_R0_clk),
    .R0_data(mem_127_1_R0_data),
    .R0_en(mem_127_1_R0_en),
    .W0_addr(mem_127_1_W0_addr),
    .W0_clk(mem_127_1_W0_clk),
    .W0_data(mem_127_1_W0_data),
    .W0_en(mem_127_1_W0_en),
    .W0_mask(mem_127_1_W0_mask)
  );
  split_mem_0_ext mem_127_2 (
    .R0_addr(mem_127_2_R0_addr),
    .R0_clk(mem_127_2_R0_clk),
    .R0_data(mem_127_2_R0_data),
    .R0_en(mem_127_2_R0_en),
    .W0_addr(mem_127_2_W0_addr),
    .W0_clk(mem_127_2_W0_clk),
    .W0_data(mem_127_2_W0_data),
    .W0_en(mem_127_2_W0_en),
    .W0_mask(mem_127_2_W0_mask)
  );
  split_mem_0_ext mem_127_3 (
    .R0_addr(mem_127_3_R0_addr),
    .R0_clk(mem_127_3_R0_clk),
    .R0_data(mem_127_3_R0_data),
    .R0_en(mem_127_3_R0_en),
    .W0_addr(mem_127_3_W0_addr),
    .W0_clk(mem_127_3_W0_clk),
    .W0_data(mem_127_3_W0_data),
    .W0_en(mem_127_3_W0_en),
    .W0_mask(mem_127_3_W0_mask)
  );
  split_mem_0_ext mem_127_4 (
    .R0_addr(mem_127_4_R0_addr),
    .R0_clk(mem_127_4_R0_clk),
    .R0_data(mem_127_4_R0_data),
    .R0_en(mem_127_4_R0_en),
    .W0_addr(mem_127_4_W0_addr),
    .W0_clk(mem_127_4_W0_clk),
    .W0_data(mem_127_4_W0_data),
    .W0_en(mem_127_4_W0_en),
    .W0_mask(mem_127_4_W0_mask)
  );
  split_mem_0_ext mem_127_5 (
    .R0_addr(mem_127_5_R0_addr),
    .R0_clk(mem_127_5_R0_clk),
    .R0_data(mem_127_5_R0_data),
    .R0_en(mem_127_5_R0_en),
    .W0_addr(mem_127_5_W0_addr),
    .W0_clk(mem_127_5_W0_clk),
    .W0_data(mem_127_5_W0_data),
    .W0_en(mem_127_5_W0_en),
    .W0_mask(mem_127_5_W0_mask)
  );
  split_mem_0_ext mem_127_6 (
    .R0_addr(mem_127_6_R0_addr),
    .R0_clk(mem_127_6_R0_clk),
    .R0_data(mem_127_6_R0_data),
    .R0_en(mem_127_6_R0_en),
    .W0_addr(mem_127_6_W0_addr),
    .W0_clk(mem_127_6_W0_clk),
    .W0_data(mem_127_6_W0_data),
    .W0_en(mem_127_6_W0_en),
    .W0_mask(mem_127_6_W0_mask)
  );
  split_mem_0_ext mem_127_7 (
    .R0_addr(mem_127_7_R0_addr),
    .R0_clk(mem_127_7_R0_clk),
    .R0_data(mem_127_7_R0_data),
    .R0_en(mem_127_7_R0_en),
    .W0_addr(mem_127_7_W0_addr),
    .W0_clk(mem_127_7_W0_clk),
    .W0_data(mem_127_7_W0_data),
    .W0_en(mem_127_7_W0_en),
    .W0_mask(mem_127_7_W0_mask)
  );
  split_mem_0_ext mem_128_0 (
    .R0_addr(mem_128_0_R0_addr),
    .R0_clk(mem_128_0_R0_clk),
    .R0_data(mem_128_0_R0_data),
    .R0_en(mem_128_0_R0_en),
    .W0_addr(mem_128_0_W0_addr),
    .W0_clk(mem_128_0_W0_clk),
    .W0_data(mem_128_0_W0_data),
    .W0_en(mem_128_0_W0_en),
    .W0_mask(mem_128_0_W0_mask)
  );
  split_mem_0_ext mem_128_1 (
    .R0_addr(mem_128_1_R0_addr),
    .R0_clk(mem_128_1_R0_clk),
    .R0_data(mem_128_1_R0_data),
    .R0_en(mem_128_1_R0_en),
    .W0_addr(mem_128_1_W0_addr),
    .W0_clk(mem_128_1_W0_clk),
    .W0_data(mem_128_1_W0_data),
    .W0_en(mem_128_1_W0_en),
    .W0_mask(mem_128_1_W0_mask)
  );
  split_mem_0_ext mem_128_2 (
    .R0_addr(mem_128_2_R0_addr),
    .R0_clk(mem_128_2_R0_clk),
    .R0_data(mem_128_2_R0_data),
    .R0_en(mem_128_2_R0_en),
    .W0_addr(mem_128_2_W0_addr),
    .W0_clk(mem_128_2_W0_clk),
    .W0_data(mem_128_2_W0_data),
    .W0_en(mem_128_2_W0_en),
    .W0_mask(mem_128_2_W0_mask)
  );
  split_mem_0_ext mem_128_3 (
    .R0_addr(mem_128_3_R0_addr),
    .R0_clk(mem_128_3_R0_clk),
    .R0_data(mem_128_3_R0_data),
    .R0_en(mem_128_3_R0_en),
    .W0_addr(mem_128_3_W0_addr),
    .W0_clk(mem_128_3_W0_clk),
    .W0_data(mem_128_3_W0_data),
    .W0_en(mem_128_3_W0_en),
    .W0_mask(mem_128_3_W0_mask)
  );
  split_mem_0_ext mem_128_4 (
    .R0_addr(mem_128_4_R0_addr),
    .R0_clk(mem_128_4_R0_clk),
    .R0_data(mem_128_4_R0_data),
    .R0_en(mem_128_4_R0_en),
    .W0_addr(mem_128_4_W0_addr),
    .W0_clk(mem_128_4_W0_clk),
    .W0_data(mem_128_4_W0_data),
    .W0_en(mem_128_4_W0_en),
    .W0_mask(mem_128_4_W0_mask)
  );
  split_mem_0_ext mem_128_5 (
    .R0_addr(mem_128_5_R0_addr),
    .R0_clk(mem_128_5_R0_clk),
    .R0_data(mem_128_5_R0_data),
    .R0_en(mem_128_5_R0_en),
    .W0_addr(mem_128_5_W0_addr),
    .W0_clk(mem_128_5_W0_clk),
    .W0_data(mem_128_5_W0_data),
    .W0_en(mem_128_5_W0_en),
    .W0_mask(mem_128_5_W0_mask)
  );
  split_mem_0_ext mem_128_6 (
    .R0_addr(mem_128_6_R0_addr),
    .R0_clk(mem_128_6_R0_clk),
    .R0_data(mem_128_6_R0_data),
    .R0_en(mem_128_6_R0_en),
    .W0_addr(mem_128_6_W0_addr),
    .W0_clk(mem_128_6_W0_clk),
    .W0_data(mem_128_6_W0_data),
    .W0_en(mem_128_6_W0_en),
    .W0_mask(mem_128_6_W0_mask)
  );
  split_mem_0_ext mem_128_7 (
    .R0_addr(mem_128_7_R0_addr),
    .R0_clk(mem_128_7_R0_clk),
    .R0_data(mem_128_7_R0_data),
    .R0_en(mem_128_7_R0_en),
    .W0_addr(mem_128_7_W0_addr),
    .W0_clk(mem_128_7_W0_clk),
    .W0_data(mem_128_7_W0_data),
    .W0_en(mem_128_7_W0_en),
    .W0_mask(mem_128_7_W0_mask)
  );
  split_mem_0_ext mem_129_0 (
    .R0_addr(mem_129_0_R0_addr),
    .R0_clk(mem_129_0_R0_clk),
    .R0_data(mem_129_0_R0_data),
    .R0_en(mem_129_0_R0_en),
    .W0_addr(mem_129_0_W0_addr),
    .W0_clk(mem_129_0_W0_clk),
    .W0_data(mem_129_0_W0_data),
    .W0_en(mem_129_0_W0_en),
    .W0_mask(mem_129_0_W0_mask)
  );
  split_mem_0_ext mem_129_1 (
    .R0_addr(mem_129_1_R0_addr),
    .R0_clk(mem_129_1_R0_clk),
    .R0_data(mem_129_1_R0_data),
    .R0_en(mem_129_1_R0_en),
    .W0_addr(mem_129_1_W0_addr),
    .W0_clk(mem_129_1_W0_clk),
    .W0_data(mem_129_1_W0_data),
    .W0_en(mem_129_1_W0_en),
    .W0_mask(mem_129_1_W0_mask)
  );
  split_mem_0_ext mem_129_2 (
    .R0_addr(mem_129_2_R0_addr),
    .R0_clk(mem_129_2_R0_clk),
    .R0_data(mem_129_2_R0_data),
    .R0_en(mem_129_2_R0_en),
    .W0_addr(mem_129_2_W0_addr),
    .W0_clk(mem_129_2_W0_clk),
    .W0_data(mem_129_2_W0_data),
    .W0_en(mem_129_2_W0_en),
    .W0_mask(mem_129_2_W0_mask)
  );
  split_mem_0_ext mem_129_3 (
    .R0_addr(mem_129_3_R0_addr),
    .R0_clk(mem_129_3_R0_clk),
    .R0_data(mem_129_3_R0_data),
    .R0_en(mem_129_3_R0_en),
    .W0_addr(mem_129_3_W0_addr),
    .W0_clk(mem_129_3_W0_clk),
    .W0_data(mem_129_3_W0_data),
    .W0_en(mem_129_3_W0_en),
    .W0_mask(mem_129_3_W0_mask)
  );
  split_mem_0_ext mem_129_4 (
    .R0_addr(mem_129_4_R0_addr),
    .R0_clk(mem_129_4_R0_clk),
    .R0_data(mem_129_4_R0_data),
    .R0_en(mem_129_4_R0_en),
    .W0_addr(mem_129_4_W0_addr),
    .W0_clk(mem_129_4_W0_clk),
    .W0_data(mem_129_4_W0_data),
    .W0_en(mem_129_4_W0_en),
    .W0_mask(mem_129_4_W0_mask)
  );
  split_mem_0_ext mem_129_5 (
    .R0_addr(mem_129_5_R0_addr),
    .R0_clk(mem_129_5_R0_clk),
    .R0_data(mem_129_5_R0_data),
    .R0_en(mem_129_5_R0_en),
    .W0_addr(mem_129_5_W0_addr),
    .W0_clk(mem_129_5_W0_clk),
    .W0_data(mem_129_5_W0_data),
    .W0_en(mem_129_5_W0_en),
    .W0_mask(mem_129_5_W0_mask)
  );
  split_mem_0_ext mem_129_6 (
    .R0_addr(mem_129_6_R0_addr),
    .R0_clk(mem_129_6_R0_clk),
    .R0_data(mem_129_6_R0_data),
    .R0_en(mem_129_6_R0_en),
    .W0_addr(mem_129_6_W0_addr),
    .W0_clk(mem_129_6_W0_clk),
    .W0_data(mem_129_6_W0_data),
    .W0_en(mem_129_6_W0_en),
    .W0_mask(mem_129_6_W0_mask)
  );
  split_mem_0_ext mem_129_7 (
    .R0_addr(mem_129_7_R0_addr),
    .R0_clk(mem_129_7_R0_clk),
    .R0_data(mem_129_7_R0_data),
    .R0_en(mem_129_7_R0_en),
    .W0_addr(mem_129_7_W0_addr),
    .W0_clk(mem_129_7_W0_clk),
    .W0_data(mem_129_7_W0_data),
    .W0_en(mem_129_7_W0_en),
    .W0_mask(mem_129_7_W0_mask)
  );
  split_mem_0_ext mem_130_0 (
    .R0_addr(mem_130_0_R0_addr),
    .R0_clk(mem_130_0_R0_clk),
    .R0_data(mem_130_0_R0_data),
    .R0_en(mem_130_0_R0_en),
    .W0_addr(mem_130_0_W0_addr),
    .W0_clk(mem_130_0_W0_clk),
    .W0_data(mem_130_0_W0_data),
    .W0_en(mem_130_0_W0_en),
    .W0_mask(mem_130_0_W0_mask)
  );
  split_mem_0_ext mem_130_1 (
    .R0_addr(mem_130_1_R0_addr),
    .R0_clk(mem_130_1_R0_clk),
    .R0_data(mem_130_1_R0_data),
    .R0_en(mem_130_1_R0_en),
    .W0_addr(mem_130_1_W0_addr),
    .W0_clk(mem_130_1_W0_clk),
    .W0_data(mem_130_1_W0_data),
    .W0_en(mem_130_1_W0_en),
    .W0_mask(mem_130_1_W0_mask)
  );
  split_mem_0_ext mem_130_2 (
    .R0_addr(mem_130_2_R0_addr),
    .R0_clk(mem_130_2_R0_clk),
    .R0_data(mem_130_2_R0_data),
    .R0_en(mem_130_2_R0_en),
    .W0_addr(mem_130_2_W0_addr),
    .W0_clk(mem_130_2_W0_clk),
    .W0_data(mem_130_2_W0_data),
    .W0_en(mem_130_2_W0_en),
    .W0_mask(mem_130_2_W0_mask)
  );
  split_mem_0_ext mem_130_3 (
    .R0_addr(mem_130_3_R0_addr),
    .R0_clk(mem_130_3_R0_clk),
    .R0_data(mem_130_3_R0_data),
    .R0_en(mem_130_3_R0_en),
    .W0_addr(mem_130_3_W0_addr),
    .W0_clk(mem_130_3_W0_clk),
    .W0_data(mem_130_3_W0_data),
    .W0_en(mem_130_3_W0_en),
    .W0_mask(mem_130_3_W0_mask)
  );
  split_mem_0_ext mem_130_4 (
    .R0_addr(mem_130_4_R0_addr),
    .R0_clk(mem_130_4_R0_clk),
    .R0_data(mem_130_4_R0_data),
    .R0_en(mem_130_4_R0_en),
    .W0_addr(mem_130_4_W0_addr),
    .W0_clk(mem_130_4_W0_clk),
    .W0_data(mem_130_4_W0_data),
    .W0_en(mem_130_4_W0_en),
    .W0_mask(mem_130_4_W0_mask)
  );
  split_mem_0_ext mem_130_5 (
    .R0_addr(mem_130_5_R0_addr),
    .R0_clk(mem_130_5_R0_clk),
    .R0_data(mem_130_5_R0_data),
    .R0_en(mem_130_5_R0_en),
    .W0_addr(mem_130_5_W0_addr),
    .W0_clk(mem_130_5_W0_clk),
    .W0_data(mem_130_5_W0_data),
    .W0_en(mem_130_5_W0_en),
    .W0_mask(mem_130_5_W0_mask)
  );
  split_mem_0_ext mem_130_6 (
    .R0_addr(mem_130_6_R0_addr),
    .R0_clk(mem_130_6_R0_clk),
    .R0_data(mem_130_6_R0_data),
    .R0_en(mem_130_6_R0_en),
    .W0_addr(mem_130_6_W0_addr),
    .W0_clk(mem_130_6_W0_clk),
    .W0_data(mem_130_6_W0_data),
    .W0_en(mem_130_6_W0_en),
    .W0_mask(mem_130_6_W0_mask)
  );
  split_mem_0_ext mem_130_7 (
    .R0_addr(mem_130_7_R0_addr),
    .R0_clk(mem_130_7_R0_clk),
    .R0_data(mem_130_7_R0_data),
    .R0_en(mem_130_7_R0_en),
    .W0_addr(mem_130_7_W0_addr),
    .W0_clk(mem_130_7_W0_clk),
    .W0_data(mem_130_7_W0_data),
    .W0_en(mem_130_7_W0_en),
    .W0_mask(mem_130_7_W0_mask)
  );
  split_mem_0_ext mem_131_0 (
    .R0_addr(mem_131_0_R0_addr),
    .R0_clk(mem_131_0_R0_clk),
    .R0_data(mem_131_0_R0_data),
    .R0_en(mem_131_0_R0_en),
    .W0_addr(mem_131_0_W0_addr),
    .W0_clk(mem_131_0_W0_clk),
    .W0_data(mem_131_0_W0_data),
    .W0_en(mem_131_0_W0_en),
    .W0_mask(mem_131_0_W0_mask)
  );
  split_mem_0_ext mem_131_1 (
    .R0_addr(mem_131_1_R0_addr),
    .R0_clk(mem_131_1_R0_clk),
    .R0_data(mem_131_1_R0_data),
    .R0_en(mem_131_1_R0_en),
    .W0_addr(mem_131_1_W0_addr),
    .W0_clk(mem_131_1_W0_clk),
    .W0_data(mem_131_1_W0_data),
    .W0_en(mem_131_1_W0_en),
    .W0_mask(mem_131_1_W0_mask)
  );
  split_mem_0_ext mem_131_2 (
    .R0_addr(mem_131_2_R0_addr),
    .R0_clk(mem_131_2_R0_clk),
    .R0_data(mem_131_2_R0_data),
    .R0_en(mem_131_2_R0_en),
    .W0_addr(mem_131_2_W0_addr),
    .W0_clk(mem_131_2_W0_clk),
    .W0_data(mem_131_2_W0_data),
    .W0_en(mem_131_2_W0_en),
    .W0_mask(mem_131_2_W0_mask)
  );
  split_mem_0_ext mem_131_3 (
    .R0_addr(mem_131_3_R0_addr),
    .R0_clk(mem_131_3_R0_clk),
    .R0_data(mem_131_3_R0_data),
    .R0_en(mem_131_3_R0_en),
    .W0_addr(mem_131_3_W0_addr),
    .W0_clk(mem_131_3_W0_clk),
    .W0_data(mem_131_3_W0_data),
    .W0_en(mem_131_3_W0_en),
    .W0_mask(mem_131_3_W0_mask)
  );
  split_mem_0_ext mem_131_4 (
    .R0_addr(mem_131_4_R0_addr),
    .R0_clk(mem_131_4_R0_clk),
    .R0_data(mem_131_4_R0_data),
    .R0_en(mem_131_4_R0_en),
    .W0_addr(mem_131_4_W0_addr),
    .W0_clk(mem_131_4_W0_clk),
    .W0_data(mem_131_4_W0_data),
    .W0_en(mem_131_4_W0_en),
    .W0_mask(mem_131_4_W0_mask)
  );
  split_mem_0_ext mem_131_5 (
    .R0_addr(mem_131_5_R0_addr),
    .R0_clk(mem_131_5_R0_clk),
    .R0_data(mem_131_5_R0_data),
    .R0_en(mem_131_5_R0_en),
    .W0_addr(mem_131_5_W0_addr),
    .W0_clk(mem_131_5_W0_clk),
    .W0_data(mem_131_5_W0_data),
    .W0_en(mem_131_5_W0_en),
    .W0_mask(mem_131_5_W0_mask)
  );
  split_mem_0_ext mem_131_6 (
    .R0_addr(mem_131_6_R0_addr),
    .R0_clk(mem_131_6_R0_clk),
    .R0_data(mem_131_6_R0_data),
    .R0_en(mem_131_6_R0_en),
    .W0_addr(mem_131_6_W0_addr),
    .W0_clk(mem_131_6_W0_clk),
    .W0_data(mem_131_6_W0_data),
    .W0_en(mem_131_6_W0_en),
    .W0_mask(mem_131_6_W0_mask)
  );
  split_mem_0_ext mem_131_7 (
    .R0_addr(mem_131_7_R0_addr),
    .R0_clk(mem_131_7_R0_clk),
    .R0_data(mem_131_7_R0_data),
    .R0_en(mem_131_7_R0_en),
    .W0_addr(mem_131_7_W0_addr),
    .W0_clk(mem_131_7_W0_clk),
    .W0_data(mem_131_7_W0_data),
    .W0_en(mem_131_7_W0_en),
    .W0_mask(mem_131_7_W0_mask)
  );
  split_mem_0_ext mem_132_0 (
    .R0_addr(mem_132_0_R0_addr),
    .R0_clk(mem_132_0_R0_clk),
    .R0_data(mem_132_0_R0_data),
    .R0_en(mem_132_0_R0_en),
    .W0_addr(mem_132_0_W0_addr),
    .W0_clk(mem_132_0_W0_clk),
    .W0_data(mem_132_0_W0_data),
    .W0_en(mem_132_0_W0_en),
    .W0_mask(mem_132_0_W0_mask)
  );
  split_mem_0_ext mem_132_1 (
    .R0_addr(mem_132_1_R0_addr),
    .R0_clk(mem_132_1_R0_clk),
    .R0_data(mem_132_1_R0_data),
    .R0_en(mem_132_1_R0_en),
    .W0_addr(mem_132_1_W0_addr),
    .W0_clk(mem_132_1_W0_clk),
    .W0_data(mem_132_1_W0_data),
    .W0_en(mem_132_1_W0_en),
    .W0_mask(mem_132_1_W0_mask)
  );
  split_mem_0_ext mem_132_2 (
    .R0_addr(mem_132_2_R0_addr),
    .R0_clk(mem_132_2_R0_clk),
    .R0_data(mem_132_2_R0_data),
    .R0_en(mem_132_2_R0_en),
    .W0_addr(mem_132_2_W0_addr),
    .W0_clk(mem_132_2_W0_clk),
    .W0_data(mem_132_2_W0_data),
    .W0_en(mem_132_2_W0_en),
    .W0_mask(mem_132_2_W0_mask)
  );
  split_mem_0_ext mem_132_3 (
    .R0_addr(mem_132_3_R0_addr),
    .R0_clk(mem_132_3_R0_clk),
    .R0_data(mem_132_3_R0_data),
    .R0_en(mem_132_3_R0_en),
    .W0_addr(mem_132_3_W0_addr),
    .W0_clk(mem_132_3_W0_clk),
    .W0_data(mem_132_3_W0_data),
    .W0_en(mem_132_3_W0_en),
    .W0_mask(mem_132_3_W0_mask)
  );
  split_mem_0_ext mem_132_4 (
    .R0_addr(mem_132_4_R0_addr),
    .R0_clk(mem_132_4_R0_clk),
    .R0_data(mem_132_4_R0_data),
    .R0_en(mem_132_4_R0_en),
    .W0_addr(mem_132_4_W0_addr),
    .W0_clk(mem_132_4_W0_clk),
    .W0_data(mem_132_4_W0_data),
    .W0_en(mem_132_4_W0_en),
    .W0_mask(mem_132_4_W0_mask)
  );
  split_mem_0_ext mem_132_5 (
    .R0_addr(mem_132_5_R0_addr),
    .R0_clk(mem_132_5_R0_clk),
    .R0_data(mem_132_5_R0_data),
    .R0_en(mem_132_5_R0_en),
    .W0_addr(mem_132_5_W0_addr),
    .W0_clk(mem_132_5_W0_clk),
    .W0_data(mem_132_5_W0_data),
    .W0_en(mem_132_5_W0_en),
    .W0_mask(mem_132_5_W0_mask)
  );
  split_mem_0_ext mem_132_6 (
    .R0_addr(mem_132_6_R0_addr),
    .R0_clk(mem_132_6_R0_clk),
    .R0_data(mem_132_6_R0_data),
    .R0_en(mem_132_6_R0_en),
    .W0_addr(mem_132_6_W0_addr),
    .W0_clk(mem_132_6_W0_clk),
    .W0_data(mem_132_6_W0_data),
    .W0_en(mem_132_6_W0_en),
    .W0_mask(mem_132_6_W0_mask)
  );
  split_mem_0_ext mem_132_7 (
    .R0_addr(mem_132_7_R0_addr),
    .R0_clk(mem_132_7_R0_clk),
    .R0_data(mem_132_7_R0_data),
    .R0_en(mem_132_7_R0_en),
    .W0_addr(mem_132_7_W0_addr),
    .W0_clk(mem_132_7_W0_clk),
    .W0_data(mem_132_7_W0_data),
    .W0_en(mem_132_7_W0_en),
    .W0_mask(mem_132_7_W0_mask)
  );
  split_mem_0_ext mem_133_0 (
    .R0_addr(mem_133_0_R0_addr),
    .R0_clk(mem_133_0_R0_clk),
    .R0_data(mem_133_0_R0_data),
    .R0_en(mem_133_0_R0_en),
    .W0_addr(mem_133_0_W0_addr),
    .W0_clk(mem_133_0_W0_clk),
    .W0_data(mem_133_0_W0_data),
    .W0_en(mem_133_0_W0_en),
    .W0_mask(mem_133_0_W0_mask)
  );
  split_mem_0_ext mem_133_1 (
    .R0_addr(mem_133_1_R0_addr),
    .R0_clk(mem_133_1_R0_clk),
    .R0_data(mem_133_1_R0_data),
    .R0_en(mem_133_1_R0_en),
    .W0_addr(mem_133_1_W0_addr),
    .W0_clk(mem_133_1_W0_clk),
    .W0_data(mem_133_1_W0_data),
    .W0_en(mem_133_1_W0_en),
    .W0_mask(mem_133_1_W0_mask)
  );
  split_mem_0_ext mem_133_2 (
    .R0_addr(mem_133_2_R0_addr),
    .R0_clk(mem_133_2_R0_clk),
    .R0_data(mem_133_2_R0_data),
    .R0_en(mem_133_2_R0_en),
    .W0_addr(mem_133_2_W0_addr),
    .W0_clk(mem_133_2_W0_clk),
    .W0_data(mem_133_2_W0_data),
    .W0_en(mem_133_2_W0_en),
    .W0_mask(mem_133_2_W0_mask)
  );
  split_mem_0_ext mem_133_3 (
    .R0_addr(mem_133_3_R0_addr),
    .R0_clk(mem_133_3_R0_clk),
    .R0_data(mem_133_3_R0_data),
    .R0_en(mem_133_3_R0_en),
    .W0_addr(mem_133_3_W0_addr),
    .W0_clk(mem_133_3_W0_clk),
    .W0_data(mem_133_3_W0_data),
    .W0_en(mem_133_3_W0_en),
    .W0_mask(mem_133_3_W0_mask)
  );
  split_mem_0_ext mem_133_4 (
    .R0_addr(mem_133_4_R0_addr),
    .R0_clk(mem_133_4_R0_clk),
    .R0_data(mem_133_4_R0_data),
    .R0_en(mem_133_4_R0_en),
    .W0_addr(mem_133_4_W0_addr),
    .W0_clk(mem_133_4_W0_clk),
    .W0_data(mem_133_4_W0_data),
    .W0_en(mem_133_4_W0_en),
    .W0_mask(mem_133_4_W0_mask)
  );
  split_mem_0_ext mem_133_5 (
    .R0_addr(mem_133_5_R0_addr),
    .R0_clk(mem_133_5_R0_clk),
    .R0_data(mem_133_5_R0_data),
    .R0_en(mem_133_5_R0_en),
    .W0_addr(mem_133_5_W0_addr),
    .W0_clk(mem_133_5_W0_clk),
    .W0_data(mem_133_5_W0_data),
    .W0_en(mem_133_5_W0_en),
    .W0_mask(mem_133_5_W0_mask)
  );
  split_mem_0_ext mem_133_6 (
    .R0_addr(mem_133_6_R0_addr),
    .R0_clk(mem_133_6_R0_clk),
    .R0_data(mem_133_6_R0_data),
    .R0_en(mem_133_6_R0_en),
    .W0_addr(mem_133_6_W0_addr),
    .W0_clk(mem_133_6_W0_clk),
    .W0_data(mem_133_6_W0_data),
    .W0_en(mem_133_6_W0_en),
    .W0_mask(mem_133_6_W0_mask)
  );
  split_mem_0_ext mem_133_7 (
    .R0_addr(mem_133_7_R0_addr),
    .R0_clk(mem_133_7_R0_clk),
    .R0_data(mem_133_7_R0_data),
    .R0_en(mem_133_7_R0_en),
    .W0_addr(mem_133_7_W0_addr),
    .W0_clk(mem_133_7_W0_clk),
    .W0_data(mem_133_7_W0_data),
    .W0_en(mem_133_7_W0_en),
    .W0_mask(mem_133_7_W0_mask)
  );
  split_mem_0_ext mem_134_0 (
    .R0_addr(mem_134_0_R0_addr),
    .R0_clk(mem_134_0_R0_clk),
    .R0_data(mem_134_0_R0_data),
    .R0_en(mem_134_0_R0_en),
    .W0_addr(mem_134_0_W0_addr),
    .W0_clk(mem_134_0_W0_clk),
    .W0_data(mem_134_0_W0_data),
    .W0_en(mem_134_0_W0_en),
    .W0_mask(mem_134_0_W0_mask)
  );
  split_mem_0_ext mem_134_1 (
    .R0_addr(mem_134_1_R0_addr),
    .R0_clk(mem_134_1_R0_clk),
    .R0_data(mem_134_1_R0_data),
    .R0_en(mem_134_1_R0_en),
    .W0_addr(mem_134_1_W0_addr),
    .W0_clk(mem_134_1_W0_clk),
    .W0_data(mem_134_1_W0_data),
    .W0_en(mem_134_1_W0_en),
    .W0_mask(mem_134_1_W0_mask)
  );
  split_mem_0_ext mem_134_2 (
    .R0_addr(mem_134_2_R0_addr),
    .R0_clk(mem_134_2_R0_clk),
    .R0_data(mem_134_2_R0_data),
    .R0_en(mem_134_2_R0_en),
    .W0_addr(mem_134_2_W0_addr),
    .W0_clk(mem_134_2_W0_clk),
    .W0_data(mem_134_2_W0_data),
    .W0_en(mem_134_2_W0_en),
    .W0_mask(mem_134_2_W0_mask)
  );
  split_mem_0_ext mem_134_3 (
    .R0_addr(mem_134_3_R0_addr),
    .R0_clk(mem_134_3_R0_clk),
    .R0_data(mem_134_3_R0_data),
    .R0_en(mem_134_3_R0_en),
    .W0_addr(mem_134_3_W0_addr),
    .W0_clk(mem_134_3_W0_clk),
    .W0_data(mem_134_3_W0_data),
    .W0_en(mem_134_3_W0_en),
    .W0_mask(mem_134_3_W0_mask)
  );
  split_mem_0_ext mem_134_4 (
    .R0_addr(mem_134_4_R0_addr),
    .R0_clk(mem_134_4_R0_clk),
    .R0_data(mem_134_4_R0_data),
    .R0_en(mem_134_4_R0_en),
    .W0_addr(mem_134_4_W0_addr),
    .W0_clk(mem_134_4_W0_clk),
    .W0_data(mem_134_4_W0_data),
    .W0_en(mem_134_4_W0_en),
    .W0_mask(mem_134_4_W0_mask)
  );
  split_mem_0_ext mem_134_5 (
    .R0_addr(mem_134_5_R0_addr),
    .R0_clk(mem_134_5_R0_clk),
    .R0_data(mem_134_5_R0_data),
    .R0_en(mem_134_5_R0_en),
    .W0_addr(mem_134_5_W0_addr),
    .W0_clk(mem_134_5_W0_clk),
    .W0_data(mem_134_5_W0_data),
    .W0_en(mem_134_5_W0_en),
    .W0_mask(mem_134_5_W0_mask)
  );
  split_mem_0_ext mem_134_6 (
    .R0_addr(mem_134_6_R0_addr),
    .R0_clk(mem_134_6_R0_clk),
    .R0_data(mem_134_6_R0_data),
    .R0_en(mem_134_6_R0_en),
    .W0_addr(mem_134_6_W0_addr),
    .W0_clk(mem_134_6_W0_clk),
    .W0_data(mem_134_6_W0_data),
    .W0_en(mem_134_6_W0_en),
    .W0_mask(mem_134_6_W0_mask)
  );
  split_mem_0_ext mem_134_7 (
    .R0_addr(mem_134_7_R0_addr),
    .R0_clk(mem_134_7_R0_clk),
    .R0_data(mem_134_7_R0_data),
    .R0_en(mem_134_7_R0_en),
    .W0_addr(mem_134_7_W0_addr),
    .W0_clk(mem_134_7_W0_clk),
    .W0_data(mem_134_7_W0_data),
    .W0_en(mem_134_7_W0_en),
    .W0_mask(mem_134_7_W0_mask)
  );
  split_mem_0_ext mem_135_0 (
    .R0_addr(mem_135_0_R0_addr),
    .R0_clk(mem_135_0_R0_clk),
    .R0_data(mem_135_0_R0_data),
    .R0_en(mem_135_0_R0_en),
    .W0_addr(mem_135_0_W0_addr),
    .W0_clk(mem_135_0_W0_clk),
    .W0_data(mem_135_0_W0_data),
    .W0_en(mem_135_0_W0_en),
    .W0_mask(mem_135_0_W0_mask)
  );
  split_mem_0_ext mem_135_1 (
    .R0_addr(mem_135_1_R0_addr),
    .R0_clk(mem_135_1_R0_clk),
    .R0_data(mem_135_1_R0_data),
    .R0_en(mem_135_1_R0_en),
    .W0_addr(mem_135_1_W0_addr),
    .W0_clk(mem_135_1_W0_clk),
    .W0_data(mem_135_1_W0_data),
    .W0_en(mem_135_1_W0_en),
    .W0_mask(mem_135_1_W0_mask)
  );
  split_mem_0_ext mem_135_2 (
    .R0_addr(mem_135_2_R0_addr),
    .R0_clk(mem_135_2_R0_clk),
    .R0_data(mem_135_2_R0_data),
    .R0_en(mem_135_2_R0_en),
    .W0_addr(mem_135_2_W0_addr),
    .W0_clk(mem_135_2_W0_clk),
    .W0_data(mem_135_2_W0_data),
    .W0_en(mem_135_2_W0_en),
    .W0_mask(mem_135_2_W0_mask)
  );
  split_mem_0_ext mem_135_3 (
    .R0_addr(mem_135_3_R0_addr),
    .R0_clk(mem_135_3_R0_clk),
    .R0_data(mem_135_3_R0_data),
    .R0_en(mem_135_3_R0_en),
    .W0_addr(mem_135_3_W0_addr),
    .W0_clk(mem_135_3_W0_clk),
    .W0_data(mem_135_3_W0_data),
    .W0_en(mem_135_3_W0_en),
    .W0_mask(mem_135_3_W0_mask)
  );
  split_mem_0_ext mem_135_4 (
    .R0_addr(mem_135_4_R0_addr),
    .R0_clk(mem_135_4_R0_clk),
    .R0_data(mem_135_4_R0_data),
    .R0_en(mem_135_4_R0_en),
    .W0_addr(mem_135_4_W0_addr),
    .W0_clk(mem_135_4_W0_clk),
    .W0_data(mem_135_4_W0_data),
    .W0_en(mem_135_4_W0_en),
    .W0_mask(mem_135_4_W0_mask)
  );
  split_mem_0_ext mem_135_5 (
    .R0_addr(mem_135_5_R0_addr),
    .R0_clk(mem_135_5_R0_clk),
    .R0_data(mem_135_5_R0_data),
    .R0_en(mem_135_5_R0_en),
    .W0_addr(mem_135_5_W0_addr),
    .W0_clk(mem_135_5_W0_clk),
    .W0_data(mem_135_5_W0_data),
    .W0_en(mem_135_5_W0_en),
    .W0_mask(mem_135_5_W0_mask)
  );
  split_mem_0_ext mem_135_6 (
    .R0_addr(mem_135_6_R0_addr),
    .R0_clk(mem_135_6_R0_clk),
    .R0_data(mem_135_6_R0_data),
    .R0_en(mem_135_6_R0_en),
    .W0_addr(mem_135_6_W0_addr),
    .W0_clk(mem_135_6_W0_clk),
    .W0_data(mem_135_6_W0_data),
    .W0_en(mem_135_6_W0_en),
    .W0_mask(mem_135_6_W0_mask)
  );
  split_mem_0_ext mem_135_7 (
    .R0_addr(mem_135_7_R0_addr),
    .R0_clk(mem_135_7_R0_clk),
    .R0_data(mem_135_7_R0_data),
    .R0_en(mem_135_7_R0_en),
    .W0_addr(mem_135_7_W0_addr),
    .W0_clk(mem_135_7_W0_clk),
    .W0_data(mem_135_7_W0_data),
    .W0_en(mem_135_7_W0_en),
    .W0_mask(mem_135_7_W0_mask)
  );
  split_mem_0_ext mem_136_0 (
    .R0_addr(mem_136_0_R0_addr),
    .R0_clk(mem_136_0_R0_clk),
    .R0_data(mem_136_0_R0_data),
    .R0_en(mem_136_0_R0_en),
    .W0_addr(mem_136_0_W0_addr),
    .W0_clk(mem_136_0_W0_clk),
    .W0_data(mem_136_0_W0_data),
    .W0_en(mem_136_0_W0_en),
    .W0_mask(mem_136_0_W0_mask)
  );
  split_mem_0_ext mem_136_1 (
    .R0_addr(mem_136_1_R0_addr),
    .R0_clk(mem_136_1_R0_clk),
    .R0_data(mem_136_1_R0_data),
    .R0_en(mem_136_1_R0_en),
    .W0_addr(mem_136_1_W0_addr),
    .W0_clk(mem_136_1_W0_clk),
    .W0_data(mem_136_1_W0_data),
    .W0_en(mem_136_1_W0_en),
    .W0_mask(mem_136_1_W0_mask)
  );
  split_mem_0_ext mem_136_2 (
    .R0_addr(mem_136_2_R0_addr),
    .R0_clk(mem_136_2_R0_clk),
    .R0_data(mem_136_2_R0_data),
    .R0_en(mem_136_2_R0_en),
    .W0_addr(mem_136_2_W0_addr),
    .W0_clk(mem_136_2_W0_clk),
    .W0_data(mem_136_2_W0_data),
    .W0_en(mem_136_2_W0_en),
    .W0_mask(mem_136_2_W0_mask)
  );
  split_mem_0_ext mem_136_3 (
    .R0_addr(mem_136_3_R0_addr),
    .R0_clk(mem_136_3_R0_clk),
    .R0_data(mem_136_3_R0_data),
    .R0_en(mem_136_3_R0_en),
    .W0_addr(mem_136_3_W0_addr),
    .W0_clk(mem_136_3_W0_clk),
    .W0_data(mem_136_3_W0_data),
    .W0_en(mem_136_3_W0_en),
    .W0_mask(mem_136_3_W0_mask)
  );
  split_mem_0_ext mem_136_4 (
    .R0_addr(mem_136_4_R0_addr),
    .R0_clk(mem_136_4_R0_clk),
    .R0_data(mem_136_4_R0_data),
    .R0_en(mem_136_4_R0_en),
    .W0_addr(mem_136_4_W0_addr),
    .W0_clk(mem_136_4_W0_clk),
    .W0_data(mem_136_4_W0_data),
    .W0_en(mem_136_4_W0_en),
    .W0_mask(mem_136_4_W0_mask)
  );
  split_mem_0_ext mem_136_5 (
    .R0_addr(mem_136_5_R0_addr),
    .R0_clk(mem_136_5_R0_clk),
    .R0_data(mem_136_5_R0_data),
    .R0_en(mem_136_5_R0_en),
    .W0_addr(mem_136_5_W0_addr),
    .W0_clk(mem_136_5_W0_clk),
    .W0_data(mem_136_5_W0_data),
    .W0_en(mem_136_5_W0_en),
    .W0_mask(mem_136_5_W0_mask)
  );
  split_mem_0_ext mem_136_6 (
    .R0_addr(mem_136_6_R0_addr),
    .R0_clk(mem_136_6_R0_clk),
    .R0_data(mem_136_6_R0_data),
    .R0_en(mem_136_6_R0_en),
    .W0_addr(mem_136_6_W0_addr),
    .W0_clk(mem_136_6_W0_clk),
    .W0_data(mem_136_6_W0_data),
    .W0_en(mem_136_6_W0_en),
    .W0_mask(mem_136_6_W0_mask)
  );
  split_mem_0_ext mem_136_7 (
    .R0_addr(mem_136_7_R0_addr),
    .R0_clk(mem_136_7_R0_clk),
    .R0_data(mem_136_7_R0_data),
    .R0_en(mem_136_7_R0_en),
    .W0_addr(mem_136_7_W0_addr),
    .W0_clk(mem_136_7_W0_clk),
    .W0_data(mem_136_7_W0_data),
    .W0_en(mem_136_7_W0_en),
    .W0_mask(mem_136_7_W0_mask)
  );
  split_mem_0_ext mem_137_0 (
    .R0_addr(mem_137_0_R0_addr),
    .R0_clk(mem_137_0_R0_clk),
    .R0_data(mem_137_0_R0_data),
    .R0_en(mem_137_0_R0_en),
    .W0_addr(mem_137_0_W0_addr),
    .W0_clk(mem_137_0_W0_clk),
    .W0_data(mem_137_0_W0_data),
    .W0_en(mem_137_0_W0_en),
    .W0_mask(mem_137_0_W0_mask)
  );
  split_mem_0_ext mem_137_1 (
    .R0_addr(mem_137_1_R0_addr),
    .R0_clk(mem_137_1_R0_clk),
    .R0_data(mem_137_1_R0_data),
    .R0_en(mem_137_1_R0_en),
    .W0_addr(mem_137_1_W0_addr),
    .W0_clk(mem_137_1_W0_clk),
    .W0_data(mem_137_1_W0_data),
    .W0_en(mem_137_1_W0_en),
    .W0_mask(mem_137_1_W0_mask)
  );
  split_mem_0_ext mem_137_2 (
    .R0_addr(mem_137_2_R0_addr),
    .R0_clk(mem_137_2_R0_clk),
    .R0_data(mem_137_2_R0_data),
    .R0_en(mem_137_2_R0_en),
    .W0_addr(mem_137_2_W0_addr),
    .W0_clk(mem_137_2_W0_clk),
    .W0_data(mem_137_2_W0_data),
    .W0_en(mem_137_2_W0_en),
    .W0_mask(mem_137_2_W0_mask)
  );
  split_mem_0_ext mem_137_3 (
    .R0_addr(mem_137_3_R0_addr),
    .R0_clk(mem_137_3_R0_clk),
    .R0_data(mem_137_3_R0_data),
    .R0_en(mem_137_3_R0_en),
    .W0_addr(mem_137_3_W0_addr),
    .W0_clk(mem_137_3_W0_clk),
    .W0_data(mem_137_3_W0_data),
    .W0_en(mem_137_3_W0_en),
    .W0_mask(mem_137_3_W0_mask)
  );
  split_mem_0_ext mem_137_4 (
    .R0_addr(mem_137_4_R0_addr),
    .R0_clk(mem_137_4_R0_clk),
    .R0_data(mem_137_4_R0_data),
    .R0_en(mem_137_4_R0_en),
    .W0_addr(mem_137_4_W0_addr),
    .W0_clk(mem_137_4_W0_clk),
    .W0_data(mem_137_4_W0_data),
    .W0_en(mem_137_4_W0_en),
    .W0_mask(mem_137_4_W0_mask)
  );
  split_mem_0_ext mem_137_5 (
    .R0_addr(mem_137_5_R0_addr),
    .R0_clk(mem_137_5_R0_clk),
    .R0_data(mem_137_5_R0_data),
    .R0_en(mem_137_5_R0_en),
    .W0_addr(mem_137_5_W0_addr),
    .W0_clk(mem_137_5_W0_clk),
    .W0_data(mem_137_5_W0_data),
    .W0_en(mem_137_5_W0_en),
    .W0_mask(mem_137_5_W0_mask)
  );
  split_mem_0_ext mem_137_6 (
    .R0_addr(mem_137_6_R0_addr),
    .R0_clk(mem_137_6_R0_clk),
    .R0_data(mem_137_6_R0_data),
    .R0_en(mem_137_6_R0_en),
    .W0_addr(mem_137_6_W0_addr),
    .W0_clk(mem_137_6_W0_clk),
    .W0_data(mem_137_6_W0_data),
    .W0_en(mem_137_6_W0_en),
    .W0_mask(mem_137_6_W0_mask)
  );
  split_mem_0_ext mem_137_7 (
    .R0_addr(mem_137_7_R0_addr),
    .R0_clk(mem_137_7_R0_clk),
    .R0_data(mem_137_7_R0_data),
    .R0_en(mem_137_7_R0_en),
    .W0_addr(mem_137_7_W0_addr),
    .W0_clk(mem_137_7_W0_clk),
    .W0_data(mem_137_7_W0_data),
    .W0_en(mem_137_7_W0_en),
    .W0_mask(mem_137_7_W0_mask)
  );
  split_mem_0_ext mem_138_0 (
    .R0_addr(mem_138_0_R0_addr),
    .R0_clk(mem_138_0_R0_clk),
    .R0_data(mem_138_0_R0_data),
    .R0_en(mem_138_0_R0_en),
    .W0_addr(mem_138_0_W0_addr),
    .W0_clk(mem_138_0_W0_clk),
    .W0_data(mem_138_0_W0_data),
    .W0_en(mem_138_0_W0_en),
    .W0_mask(mem_138_0_W0_mask)
  );
  split_mem_0_ext mem_138_1 (
    .R0_addr(mem_138_1_R0_addr),
    .R0_clk(mem_138_1_R0_clk),
    .R0_data(mem_138_1_R0_data),
    .R0_en(mem_138_1_R0_en),
    .W0_addr(mem_138_1_W0_addr),
    .W0_clk(mem_138_1_W0_clk),
    .W0_data(mem_138_1_W0_data),
    .W0_en(mem_138_1_W0_en),
    .W0_mask(mem_138_1_W0_mask)
  );
  split_mem_0_ext mem_138_2 (
    .R0_addr(mem_138_2_R0_addr),
    .R0_clk(mem_138_2_R0_clk),
    .R0_data(mem_138_2_R0_data),
    .R0_en(mem_138_2_R0_en),
    .W0_addr(mem_138_2_W0_addr),
    .W0_clk(mem_138_2_W0_clk),
    .W0_data(mem_138_2_W0_data),
    .W0_en(mem_138_2_W0_en),
    .W0_mask(mem_138_2_W0_mask)
  );
  split_mem_0_ext mem_138_3 (
    .R0_addr(mem_138_3_R0_addr),
    .R0_clk(mem_138_3_R0_clk),
    .R0_data(mem_138_3_R0_data),
    .R0_en(mem_138_3_R0_en),
    .W0_addr(mem_138_3_W0_addr),
    .W0_clk(mem_138_3_W0_clk),
    .W0_data(mem_138_3_W0_data),
    .W0_en(mem_138_3_W0_en),
    .W0_mask(mem_138_3_W0_mask)
  );
  split_mem_0_ext mem_138_4 (
    .R0_addr(mem_138_4_R0_addr),
    .R0_clk(mem_138_4_R0_clk),
    .R0_data(mem_138_4_R0_data),
    .R0_en(mem_138_4_R0_en),
    .W0_addr(mem_138_4_W0_addr),
    .W0_clk(mem_138_4_W0_clk),
    .W0_data(mem_138_4_W0_data),
    .W0_en(mem_138_4_W0_en),
    .W0_mask(mem_138_4_W0_mask)
  );
  split_mem_0_ext mem_138_5 (
    .R0_addr(mem_138_5_R0_addr),
    .R0_clk(mem_138_5_R0_clk),
    .R0_data(mem_138_5_R0_data),
    .R0_en(mem_138_5_R0_en),
    .W0_addr(mem_138_5_W0_addr),
    .W0_clk(mem_138_5_W0_clk),
    .W0_data(mem_138_5_W0_data),
    .W0_en(mem_138_5_W0_en),
    .W0_mask(mem_138_5_W0_mask)
  );
  split_mem_0_ext mem_138_6 (
    .R0_addr(mem_138_6_R0_addr),
    .R0_clk(mem_138_6_R0_clk),
    .R0_data(mem_138_6_R0_data),
    .R0_en(mem_138_6_R0_en),
    .W0_addr(mem_138_6_W0_addr),
    .W0_clk(mem_138_6_W0_clk),
    .W0_data(mem_138_6_W0_data),
    .W0_en(mem_138_6_W0_en),
    .W0_mask(mem_138_6_W0_mask)
  );
  split_mem_0_ext mem_138_7 (
    .R0_addr(mem_138_7_R0_addr),
    .R0_clk(mem_138_7_R0_clk),
    .R0_data(mem_138_7_R0_data),
    .R0_en(mem_138_7_R0_en),
    .W0_addr(mem_138_7_W0_addr),
    .W0_clk(mem_138_7_W0_clk),
    .W0_data(mem_138_7_W0_data),
    .W0_en(mem_138_7_W0_en),
    .W0_mask(mem_138_7_W0_mask)
  );
  split_mem_0_ext mem_139_0 (
    .R0_addr(mem_139_0_R0_addr),
    .R0_clk(mem_139_0_R0_clk),
    .R0_data(mem_139_0_R0_data),
    .R0_en(mem_139_0_R0_en),
    .W0_addr(mem_139_0_W0_addr),
    .W0_clk(mem_139_0_W0_clk),
    .W0_data(mem_139_0_W0_data),
    .W0_en(mem_139_0_W0_en),
    .W0_mask(mem_139_0_W0_mask)
  );
  split_mem_0_ext mem_139_1 (
    .R0_addr(mem_139_1_R0_addr),
    .R0_clk(mem_139_1_R0_clk),
    .R0_data(mem_139_1_R0_data),
    .R0_en(mem_139_1_R0_en),
    .W0_addr(mem_139_1_W0_addr),
    .W0_clk(mem_139_1_W0_clk),
    .W0_data(mem_139_1_W0_data),
    .W0_en(mem_139_1_W0_en),
    .W0_mask(mem_139_1_W0_mask)
  );
  split_mem_0_ext mem_139_2 (
    .R0_addr(mem_139_2_R0_addr),
    .R0_clk(mem_139_2_R0_clk),
    .R0_data(mem_139_2_R0_data),
    .R0_en(mem_139_2_R0_en),
    .W0_addr(mem_139_2_W0_addr),
    .W0_clk(mem_139_2_W0_clk),
    .W0_data(mem_139_2_W0_data),
    .W0_en(mem_139_2_W0_en),
    .W0_mask(mem_139_2_W0_mask)
  );
  split_mem_0_ext mem_139_3 (
    .R0_addr(mem_139_3_R0_addr),
    .R0_clk(mem_139_3_R0_clk),
    .R0_data(mem_139_3_R0_data),
    .R0_en(mem_139_3_R0_en),
    .W0_addr(mem_139_3_W0_addr),
    .W0_clk(mem_139_3_W0_clk),
    .W0_data(mem_139_3_W0_data),
    .W0_en(mem_139_3_W0_en),
    .W0_mask(mem_139_3_W0_mask)
  );
  split_mem_0_ext mem_139_4 (
    .R0_addr(mem_139_4_R0_addr),
    .R0_clk(mem_139_4_R0_clk),
    .R0_data(mem_139_4_R0_data),
    .R0_en(mem_139_4_R0_en),
    .W0_addr(mem_139_4_W0_addr),
    .W0_clk(mem_139_4_W0_clk),
    .W0_data(mem_139_4_W0_data),
    .W0_en(mem_139_4_W0_en),
    .W0_mask(mem_139_4_W0_mask)
  );
  split_mem_0_ext mem_139_5 (
    .R0_addr(mem_139_5_R0_addr),
    .R0_clk(mem_139_5_R0_clk),
    .R0_data(mem_139_5_R0_data),
    .R0_en(mem_139_5_R0_en),
    .W0_addr(mem_139_5_W0_addr),
    .W0_clk(mem_139_5_W0_clk),
    .W0_data(mem_139_5_W0_data),
    .W0_en(mem_139_5_W0_en),
    .W0_mask(mem_139_5_W0_mask)
  );
  split_mem_0_ext mem_139_6 (
    .R0_addr(mem_139_6_R0_addr),
    .R0_clk(mem_139_6_R0_clk),
    .R0_data(mem_139_6_R0_data),
    .R0_en(mem_139_6_R0_en),
    .W0_addr(mem_139_6_W0_addr),
    .W0_clk(mem_139_6_W0_clk),
    .W0_data(mem_139_6_W0_data),
    .W0_en(mem_139_6_W0_en),
    .W0_mask(mem_139_6_W0_mask)
  );
  split_mem_0_ext mem_139_7 (
    .R0_addr(mem_139_7_R0_addr),
    .R0_clk(mem_139_7_R0_clk),
    .R0_data(mem_139_7_R0_data),
    .R0_en(mem_139_7_R0_en),
    .W0_addr(mem_139_7_W0_addr),
    .W0_clk(mem_139_7_W0_clk),
    .W0_data(mem_139_7_W0_data),
    .W0_en(mem_139_7_W0_en),
    .W0_mask(mem_139_7_W0_mask)
  );
  split_mem_0_ext mem_140_0 (
    .R0_addr(mem_140_0_R0_addr),
    .R0_clk(mem_140_0_R0_clk),
    .R0_data(mem_140_0_R0_data),
    .R0_en(mem_140_0_R0_en),
    .W0_addr(mem_140_0_W0_addr),
    .W0_clk(mem_140_0_W0_clk),
    .W0_data(mem_140_0_W0_data),
    .W0_en(mem_140_0_W0_en),
    .W0_mask(mem_140_0_W0_mask)
  );
  split_mem_0_ext mem_140_1 (
    .R0_addr(mem_140_1_R0_addr),
    .R0_clk(mem_140_1_R0_clk),
    .R0_data(mem_140_1_R0_data),
    .R0_en(mem_140_1_R0_en),
    .W0_addr(mem_140_1_W0_addr),
    .W0_clk(mem_140_1_W0_clk),
    .W0_data(mem_140_1_W0_data),
    .W0_en(mem_140_1_W0_en),
    .W0_mask(mem_140_1_W0_mask)
  );
  split_mem_0_ext mem_140_2 (
    .R0_addr(mem_140_2_R0_addr),
    .R0_clk(mem_140_2_R0_clk),
    .R0_data(mem_140_2_R0_data),
    .R0_en(mem_140_2_R0_en),
    .W0_addr(mem_140_2_W0_addr),
    .W0_clk(mem_140_2_W0_clk),
    .W0_data(mem_140_2_W0_data),
    .W0_en(mem_140_2_W0_en),
    .W0_mask(mem_140_2_W0_mask)
  );
  split_mem_0_ext mem_140_3 (
    .R0_addr(mem_140_3_R0_addr),
    .R0_clk(mem_140_3_R0_clk),
    .R0_data(mem_140_3_R0_data),
    .R0_en(mem_140_3_R0_en),
    .W0_addr(mem_140_3_W0_addr),
    .W0_clk(mem_140_3_W0_clk),
    .W0_data(mem_140_3_W0_data),
    .W0_en(mem_140_3_W0_en),
    .W0_mask(mem_140_3_W0_mask)
  );
  split_mem_0_ext mem_140_4 (
    .R0_addr(mem_140_4_R0_addr),
    .R0_clk(mem_140_4_R0_clk),
    .R0_data(mem_140_4_R0_data),
    .R0_en(mem_140_4_R0_en),
    .W0_addr(mem_140_4_W0_addr),
    .W0_clk(mem_140_4_W0_clk),
    .W0_data(mem_140_4_W0_data),
    .W0_en(mem_140_4_W0_en),
    .W0_mask(mem_140_4_W0_mask)
  );
  split_mem_0_ext mem_140_5 (
    .R0_addr(mem_140_5_R0_addr),
    .R0_clk(mem_140_5_R0_clk),
    .R0_data(mem_140_5_R0_data),
    .R0_en(mem_140_5_R0_en),
    .W0_addr(mem_140_5_W0_addr),
    .W0_clk(mem_140_5_W0_clk),
    .W0_data(mem_140_5_W0_data),
    .W0_en(mem_140_5_W0_en),
    .W0_mask(mem_140_5_W0_mask)
  );
  split_mem_0_ext mem_140_6 (
    .R0_addr(mem_140_6_R0_addr),
    .R0_clk(mem_140_6_R0_clk),
    .R0_data(mem_140_6_R0_data),
    .R0_en(mem_140_6_R0_en),
    .W0_addr(mem_140_6_W0_addr),
    .W0_clk(mem_140_6_W0_clk),
    .W0_data(mem_140_6_W0_data),
    .W0_en(mem_140_6_W0_en),
    .W0_mask(mem_140_6_W0_mask)
  );
  split_mem_0_ext mem_140_7 (
    .R0_addr(mem_140_7_R0_addr),
    .R0_clk(mem_140_7_R0_clk),
    .R0_data(mem_140_7_R0_data),
    .R0_en(mem_140_7_R0_en),
    .W0_addr(mem_140_7_W0_addr),
    .W0_clk(mem_140_7_W0_clk),
    .W0_data(mem_140_7_W0_data),
    .W0_en(mem_140_7_W0_en),
    .W0_mask(mem_140_7_W0_mask)
  );
  split_mem_0_ext mem_141_0 (
    .R0_addr(mem_141_0_R0_addr),
    .R0_clk(mem_141_0_R0_clk),
    .R0_data(mem_141_0_R0_data),
    .R0_en(mem_141_0_R0_en),
    .W0_addr(mem_141_0_W0_addr),
    .W0_clk(mem_141_0_W0_clk),
    .W0_data(mem_141_0_W0_data),
    .W0_en(mem_141_0_W0_en),
    .W0_mask(mem_141_0_W0_mask)
  );
  split_mem_0_ext mem_141_1 (
    .R0_addr(mem_141_1_R0_addr),
    .R0_clk(mem_141_1_R0_clk),
    .R0_data(mem_141_1_R0_data),
    .R0_en(mem_141_1_R0_en),
    .W0_addr(mem_141_1_W0_addr),
    .W0_clk(mem_141_1_W0_clk),
    .W0_data(mem_141_1_W0_data),
    .W0_en(mem_141_1_W0_en),
    .W0_mask(mem_141_1_W0_mask)
  );
  split_mem_0_ext mem_141_2 (
    .R0_addr(mem_141_2_R0_addr),
    .R0_clk(mem_141_2_R0_clk),
    .R0_data(mem_141_2_R0_data),
    .R0_en(mem_141_2_R0_en),
    .W0_addr(mem_141_2_W0_addr),
    .W0_clk(mem_141_2_W0_clk),
    .W0_data(mem_141_2_W0_data),
    .W0_en(mem_141_2_W0_en),
    .W0_mask(mem_141_2_W0_mask)
  );
  split_mem_0_ext mem_141_3 (
    .R0_addr(mem_141_3_R0_addr),
    .R0_clk(mem_141_3_R0_clk),
    .R0_data(mem_141_3_R0_data),
    .R0_en(mem_141_3_R0_en),
    .W0_addr(mem_141_3_W0_addr),
    .W0_clk(mem_141_3_W0_clk),
    .W0_data(mem_141_3_W0_data),
    .W0_en(mem_141_3_W0_en),
    .W0_mask(mem_141_3_W0_mask)
  );
  split_mem_0_ext mem_141_4 (
    .R0_addr(mem_141_4_R0_addr),
    .R0_clk(mem_141_4_R0_clk),
    .R0_data(mem_141_4_R0_data),
    .R0_en(mem_141_4_R0_en),
    .W0_addr(mem_141_4_W0_addr),
    .W0_clk(mem_141_4_W0_clk),
    .W0_data(mem_141_4_W0_data),
    .W0_en(mem_141_4_W0_en),
    .W0_mask(mem_141_4_W0_mask)
  );
  split_mem_0_ext mem_141_5 (
    .R0_addr(mem_141_5_R0_addr),
    .R0_clk(mem_141_5_R0_clk),
    .R0_data(mem_141_5_R0_data),
    .R0_en(mem_141_5_R0_en),
    .W0_addr(mem_141_5_W0_addr),
    .W0_clk(mem_141_5_W0_clk),
    .W0_data(mem_141_5_W0_data),
    .W0_en(mem_141_5_W0_en),
    .W0_mask(mem_141_5_W0_mask)
  );
  split_mem_0_ext mem_141_6 (
    .R0_addr(mem_141_6_R0_addr),
    .R0_clk(mem_141_6_R0_clk),
    .R0_data(mem_141_6_R0_data),
    .R0_en(mem_141_6_R0_en),
    .W0_addr(mem_141_6_W0_addr),
    .W0_clk(mem_141_6_W0_clk),
    .W0_data(mem_141_6_W0_data),
    .W0_en(mem_141_6_W0_en),
    .W0_mask(mem_141_6_W0_mask)
  );
  split_mem_0_ext mem_141_7 (
    .R0_addr(mem_141_7_R0_addr),
    .R0_clk(mem_141_7_R0_clk),
    .R0_data(mem_141_7_R0_data),
    .R0_en(mem_141_7_R0_en),
    .W0_addr(mem_141_7_W0_addr),
    .W0_clk(mem_141_7_W0_clk),
    .W0_data(mem_141_7_W0_data),
    .W0_en(mem_141_7_W0_en),
    .W0_mask(mem_141_7_W0_mask)
  );
  split_mem_0_ext mem_142_0 (
    .R0_addr(mem_142_0_R0_addr),
    .R0_clk(mem_142_0_R0_clk),
    .R0_data(mem_142_0_R0_data),
    .R0_en(mem_142_0_R0_en),
    .W0_addr(mem_142_0_W0_addr),
    .W0_clk(mem_142_0_W0_clk),
    .W0_data(mem_142_0_W0_data),
    .W0_en(mem_142_0_W0_en),
    .W0_mask(mem_142_0_W0_mask)
  );
  split_mem_0_ext mem_142_1 (
    .R0_addr(mem_142_1_R0_addr),
    .R0_clk(mem_142_1_R0_clk),
    .R0_data(mem_142_1_R0_data),
    .R0_en(mem_142_1_R0_en),
    .W0_addr(mem_142_1_W0_addr),
    .W0_clk(mem_142_1_W0_clk),
    .W0_data(mem_142_1_W0_data),
    .W0_en(mem_142_1_W0_en),
    .W0_mask(mem_142_1_W0_mask)
  );
  split_mem_0_ext mem_142_2 (
    .R0_addr(mem_142_2_R0_addr),
    .R0_clk(mem_142_2_R0_clk),
    .R0_data(mem_142_2_R0_data),
    .R0_en(mem_142_2_R0_en),
    .W0_addr(mem_142_2_W0_addr),
    .W0_clk(mem_142_2_W0_clk),
    .W0_data(mem_142_2_W0_data),
    .W0_en(mem_142_2_W0_en),
    .W0_mask(mem_142_2_W0_mask)
  );
  split_mem_0_ext mem_142_3 (
    .R0_addr(mem_142_3_R0_addr),
    .R0_clk(mem_142_3_R0_clk),
    .R0_data(mem_142_3_R0_data),
    .R0_en(mem_142_3_R0_en),
    .W0_addr(mem_142_3_W0_addr),
    .W0_clk(mem_142_3_W0_clk),
    .W0_data(mem_142_3_W0_data),
    .W0_en(mem_142_3_W0_en),
    .W0_mask(mem_142_3_W0_mask)
  );
  split_mem_0_ext mem_142_4 (
    .R0_addr(mem_142_4_R0_addr),
    .R0_clk(mem_142_4_R0_clk),
    .R0_data(mem_142_4_R0_data),
    .R0_en(mem_142_4_R0_en),
    .W0_addr(mem_142_4_W0_addr),
    .W0_clk(mem_142_4_W0_clk),
    .W0_data(mem_142_4_W0_data),
    .W0_en(mem_142_4_W0_en),
    .W0_mask(mem_142_4_W0_mask)
  );
  split_mem_0_ext mem_142_5 (
    .R0_addr(mem_142_5_R0_addr),
    .R0_clk(mem_142_5_R0_clk),
    .R0_data(mem_142_5_R0_data),
    .R0_en(mem_142_5_R0_en),
    .W0_addr(mem_142_5_W0_addr),
    .W0_clk(mem_142_5_W0_clk),
    .W0_data(mem_142_5_W0_data),
    .W0_en(mem_142_5_W0_en),
    .W0_mask(mem_142_5_W0_mask)
  );
  split_mem_0_ext mem_142_6 (
    .R0_addr(mem_142_6_R0_addr),
    .R0_clk(mem_142_6_R0_clk),
    .R0_data(mem_142_6_R0_data),
    .R0_en(mem_142_6_R0_en),
    .W0_addr(mem_142_6_W0_addr),
    .W0_clk(mem_142_6_W0_clk),
    .W0_data(mem_142_6_W0_data),
    .W0_en(mem_142_6_W0_en),
    .W0_mask(mem_142_6_W0_mask)
  );
  split_mem_0_ext mem_142_7 (
    .R0_addr(mem_142_7_R0_addr),
    .R0_clk(mem_142_7_R0_clk),
    .R0_data(mem_142_7_R0_data),
    .R0_en(mem_142_7_R0_en),
    .W0_addr(mem_142_7_W0_addr),
    .W0_clk(mem_142_7_W0_clk),
    .W0_data(mem_142_7_W0_data),
    .W0_en(mem_142_7_W0_en),
    .W0_mask(mem_142_7_W0_mask)
  );
  split_mem_0_ext mem_143_0 (
    .R0_addr(mem_143_0_R0_addr),
    .R0_clk(mem_143_0_R0_clk),
    .R0_data(mem_143_0_R0_data),
    .R0_en(mem_143_0_R0_en),
    .W0_addr(mem_143_0_W0_addr),
    .W0_clk(mem_143_0_W0_clk),
    .W0_data(mem_143_0_W0_data),
    .W0_en(mem_143_0_W0_en),
    .W0_mask(mem_143_0_W0_mask)
  );
  split_mem_0_ext mem_143_1 (
    .R0_addr(mem_143_1_R0_addr),
    .R0_clk(mem_143_1_R0_clk),
    .R0_data(mem_143_1_R0_data),
    .R0_en(mem_143_1_R0_en),
    .W0_addr(mem_143_1_W0_addr),
    .W0_clk(mem_143_1_W0_clk),
    .W0_data(mem_143_1_W0_data),
    .W0_en(mem_143_1_W0_en),
    .W0_mask(mem_143_1_W0_mask)
  );
  split_mem_0_ext mem_143_2 (
    .R0_addr(mem_143_2_R0_addr),
    .R0_clk(mem_143_2_R0_clk),
    .R0_data(mem_143_2_R0_data),
    .R0_en(mem_143_2_R0_en),
    .W0_addr(mem_143_2_W0_addr),
    .W0_clk(mem_143_2_W0_clk),
    .W0_data(mem_143_2_W0_data),
    .W0_en(mem_143_2_W0_en),
    .W0_mask(mem_143_2_W0_mask)
  );
  split_mem_0_ext mem_143_3 (
    .R0_addr(mem_143_3_R0_addr),
    .R0_clk(mem_143_3_R0_clk),
    .R0_data(mem_143_3_R0_data),
    .R0_en(mem_143_3_R0_en),
    .W0_addr(mem_143_3_W0_addr),
    .W0_clk(mem_143_3_W0_clk),
    .W0_data(mem_143_3_W0_data),
    .W0_en(mem_143_3_W0_en),
    .W0_mask(mem_143_3_W0_mask)
  );
  split_mem_0_ext mem_143_4 (
    .R0_addr(mem_143_4_R0_addr),
    .R0_clk(mem_143_4_R0_clk),
    .R0_data(mem_143_4_R0_data),
    .R0_en(mem_143_4_R0_en),
    .W0_addr(mem_143_4_W0_addr),
    .W0_clk(mem_143_4_W0_clk),
    .W0_data(mem_143_4_W0_data),
    .W0_en(mem_143_4_W0_en),
    .W0_mask(mem_143_4_W0_mask)
  );
  split_mem_0_ext mem_143_5 (
    .R0_addr(mem_143_5_R0_addr),
    .R0_clk(mem_143_5_R0_clk),
    .R0_data(mem_143_5_R0_data),
    .R0_en(mem_143_5_R0_en),
    .W0_addr(mem_143_5_W0_addr),
    .W0_clk(mem_143_5_W0_clk),
    .W0_data(mem_143_5_W0_data),
    .W0_en(mem_143_5_W0_en),
    .W0_mask(mem_143_5_W0_mask)
  );
  split_mem_0_ext mem_143_6 (
    .R0_addr(mem_143_6_R0_addr),
    .R0_clk(mem_143_6_R0_clk),
    .R0_data(mem_143_6_R0_data),
    .R0_en(mem_143_6_R0_en),
    .W0_addr(mem_143_6_W0_addr),
    .W0_clk(mem_143_6_W0_clk),
    .W0_data(mem_143_6_W0_data),
    .W0_en(mem_143_6_W0_en),
    .W0_mask(mem_143_6_W0_mask)
  );
  split_mem_0_ext mem_143_7 (
    .R0_addr(mem_143_7_R0_addr),
    .R0_clk(mem_143_7_R0_clk),
    .R0_data(mem_143_7_R0_data),
    .R0_en(mem_143_7_R0_en),
    .W0_addr(mem_143_7_W0_addr),
    .W0_clk(mem_143_7_W0_clk),
    .W0_data(mem_143_7_W0_data),
    .W0_en(mem_143_7_W0_en),
    .W0_mask(mem_143_7_W0_mask)
  );
  split_mem_0_ext mem_144_0 (
    .R0_addr(mem_144_0_R0_addr),
    .R0_clk(mem_144_0_R0_clk),
    .R0_data(mem_144_0_R0_data),
    .R0_en(mem_144_0_R0_en),
    .W0_addr(mem_144_0_W0_addr),
    .W0_clk(mem_144_0_W0_clk),
    .W0_data(mem_144_0_W0_data),
    .W0_en(mem_144_0_W0_en),
    .W0_mask(mem_144_0_W0_mask)
  );
  split_mem_0_ext mem_144_1 (
    .R0_addr(mem_144_1_R0_addr),
    .R0_clk(mem_144_1_R0_clk),
    .R0_data(mem_144_1_R0_data),
    .R0_en(mem_144_1_R0_en),
    .W0_addr(mem_144_1_W0_addr),
    .W0_clk(mem_144_1_W0_clk),
    .W0_data(mem_144_1_W0_data),
    .W0_en(mem_144_1_W0_en),
    .W0_mask(mem_144_1_W0_mask)
  );
  split_mem_0_ext mem_144_2 (
    .R0_addr(mem_144_2_R0_addr),
    .R0_clk(mem_144_2_R0_clk),
    .R0_data(mem_144_2_R0_data),
    .R0_en(mem_144_2_R0_en),
    .W0_addr(mem_144_2_W0_addr),
    .W0_clk(mem_144_2_W0_clk),
    .W0_data(mem_144_2_W0_data),
    .W0_en(mem_144_2_W0_en),
    .W0_mask(mem_144_2_W0_mask)
  );
  split_mem_0_ext mem_144_3 (
    .R0_addr(mem_144_3_R0_addr),
    .R0_clk(mem_144_3_R0_clk),
    .R0_data(mem_144_3_R0_data),
    .R0_en(mem_144_3_R0_en),
    .W0_addr(mem_144_3_W0_addr),
    .W0_clk(mem_144_3_W0_clk),
    .W0_data(mem_144_3_W0_data),
    .W0_en(mem_144_3_W0_en),
    .W0_mask(mem_144_3_W0_mask)
  );
  split_mem_0_ext mem_144_4 (
    .R0_addr(mem_144_4_R0_addr),
    .R0_clk(mem_144_4_R0_clk),
    .R0_data(mem_144_4_R0_data),
    .R0_en(mem_144_4_R0_en),
    .W0_addr(mem_144_4_W0_addr),
    .W0_clk(mem_144_4_W0_clk),
    .W0_data(mem_144_4_W0_data),
    .W0_en(mem_144_4_W0_en),
    .W0_mask(mem_144_4_W0_mask)
  );
  split_mem_0_ext mem_144_5 (
    .R0_addr(mem_144_5_R0_addr),
    .R0_clk(mem_144_5_R0_clk),
    .R0_data(mem_144_5_R0_data),
    .R0_en(mem_144_5_R0_en),
    .W0_addr(mem_144_5_W0_addr),
    .W0_clk(mem_144_5_W0_clk),
    .W0_data(mem_144_5_W0_data),
    .W0_en(mem_144_5_W0_en),
    .W0_mask(mem_144_5_W0_mask)
  );
  split_mem_0_ext mem_144_6 (
    .R0_addr(mem_144_6_R0_addr),
    .R0_clk(mem_144_6_R0_clk),
    .R0_data(mem_144_6_R0_data),
    .R0_en(mem_144_6_R0_en),
    .W0_addr(mem_144_6_W0_addr),
    .W0_clk(mem_144_6_W0_clk),
    .W0_data(mem_144_6_W0_data),
    .W0_en(mem_144_6_W0_en),
    .W0_mask(mem_144_6_W0_mask)
  );
  split_mem_0_ext mem_144_7 (
    .R0_addr(mem_144_7_R0_addr),
    .R0_clk(mem_144_7_R0_clk),
    .R0_data(mem_144_7_R0_data),
    .R0_en(mem_144_7_R0_en),
    .W0_addr(mem_144_7_W0_addr),
    .W0_clk(mem_144_7_W0_clk),
    .W0_data(mem_144_7_W0_data),
    .W0_en(mem_144_7_W0_en),
    .W0_mask(mem_144_7_W0_mask)
  );
  split_mem_0_ext mem_145_0 (
    .R0_addr(mem_145_0_R0_addr),
    .R0_clk(mem_145_0_R0_clk),
    .R0_data(mem_145_0_R0_data),
    .R0_en(mem_145_0_R0_en),
    .W0_addr(mem_145_0_W0_addr),
    .W0_clk(mem_145_0_W0_clk),
    .W0_data(mem_145_0_W0_data),
    .W0_en(mem_145_0_W0_en),
    .W0_mask(mem_145_0_W0_mask)
  );
  split_mem_0_ext mem_145_1 (
    .R0_addr(mem_145_1_R0_addr),
    .R0_clk(mem_145_1_R0_clk),
    .R0_data(mem_145_1_R0_data),
    .R0_en(mem_145_1_R0_en),
    .W0_addr(mem_145_1_W0_addr),
    .W0_clk(mem_145_1_W0_clk),
    .W0_data(mem_145_1_W0_data),
    .W0_en(mem_145_1_W0_en),
    .W0_mask(mem_145_1_W0_mask)
  );
  split_mem_0_ext mem_145_2 (
    .R0_addr(mem_145_2_R0_addr),
    .R0_clk(mem_145_2_R0_clk),
    .R0_data(mem_145_2_R0_data),
    .R0_en(mem_145_2_R0_en),
    .W0_addr(mem_145_2_W0_addr),
    .W0_clk(mem_145_2_W0_clk),
    .W0_data(mem_145_2_W0_data),
    .W0_en(mem_145_2_W0_en),
    .W0_mask(mem_145_2_W0_mask)
  );
  split_mem_0_ext mem_145_3 (
    .R0_addr(mem_145_3_R0_addr),
    .R0_clk(mem_145_3_R0_clk),
    .R0_data(mem_145_3_R0_data),
    .R0_en(mem_145_3_R0_en),
    .W0_addr(mem_145_3_W0_addr),
    .W0_clk(mem_145_3_W0_clk),
    .W0_data(mem_145_3_W0_data),
    .W0_en(mem_145_3_W0_en),
    .W0_mask(mem_145_3_W0_mask)
  );
  split_mem_0_ext mem_145_4 (
    .R0_addr(mem_145_4_R0_addr),
    .R0_clk(mem_145_4_R0_clk),
    .R0_data(mem_145_4_R0_data),
    .R0_en(mem_145_4_R0_en),
    .W0_addr(mem_145_4_W0_addr),
    .W0_clk(mem_145_4_W0_clk),
    .W0_data(mem_145_4_W0_data),
    .W0_en(mem_145_4_W0_en),
    .W0_mask(mem_145_4_W0_mask)
  );
  split_mem_0_ext mem_145_5 (
    .R0_addr(mem_145_5_R0_addr),
    .R0_clk(mem_145_5_R0_clk),
    .R0_data(mem_145_5_R0_data),
    .R0_en(mem_145_5_R0_en),
    .W0_addr(mem_145_5_W0_addr),
    .W0_clk(mem_145_5_W0_clk),
    .W0_data(mem_145_5_W0_data),
    .W0_en(mem_145_5_W0_en),
    .W0_mask(mem_145_5_W0_mask)
  );
  split_mem_0_ext mem_145_6 (
    .R0_addr(mem_145_6_R0_addr),
    .R0_clk(mem_145_6_R0_clk),
    .R0_data(mem_145_6_R0_data),
    .R0_en(mem_145_6_R0_en),
    .W0_addr(mem_145_6_W0_addr),
    .W0_clk(mem_145_6_W0_clk),
    .W0_data(mem_145_6_W0_data),
    .W0_en(mem_145_6_W0_en),
    .W0_mask(mem_145_6_W0_mask)
  );
  split_mem_0_ext mem_145_7 (
    .R0_addr(mem_145_7_R0_addr),
    .R0_clk(mem_145_7_R0_clk),
    .R0_data(mem_145_7_R0_data),
    .R0_en(mem_145_7_R0_en),
    .W0_addr(mem_145_7_W0_addr),
    .W0_clk(mem_145_7_W0_clk),
    .W0_data(mem_145_7_W0_data),
    .W0_en(mem_145_7_W0_en),
    .W0_mask(mem_145_7_W0_mask)
  );
  split_mem_0_ext mem_146_0 (
    .R0_addr(mem_146_0_R0_addr),
    .R0_clk(mem_146_0_R0_clk),
    .R0_data(mem_146_0_R0_data),
    .R0_en(mem_146_0_R0_en),
    .W0_addr(mem_146_0_W0_addr),
    .W0_clk(mem_146_0_W0_clk),
    .W0_data(mem_146_0_W0_data),
    .W0_en(mem_146_0_W0_en),
    .W0_mask(mem_146_0_W0_mask)
  );
  split_mem_0_ext mem_146_1 (
    .R0_addr(mem_146_1_R0_addr),
    .R0_clk(mem_146_1_R0_clk),
    .R0_data(mem_146_1_R0_data),
    .R0_en(mem_146_1_R0_en),
    .W0_addr(mem_146_1_W0_addr),
    .W0_clk(mem_146_1_W0_clk),
    .W0_data(mem_146_1_W0_data),
    .W0_en(mem_146_1_W0_en),
    .W0_mask(mem_146_1_W0_mask)
  );
  split_mem_0_ext mem_146_2 (
    .R0_addr(mem_146_2_R0_addr),
    .R0_clk(mem_146_2_R0_clk),
    .R0_data(mem_146_2_R0_data),
    .R0_en(mem_146_2_R0_en),
    .W0_addr(mem_146_2_W0_addr),
    .W0_clk(mem_146_2_W0_clk),
    .W0_data(mem_146_2_W0_data),
    .W0_en(mem_146_2_W0_en),
    .W0_mask(mem_146_2_W0_mask)
  );
  split_mem_0_ext mem_146_3 (
    .R0_addr(mem_146_3_R0_addr),
    .R0_clk(mem_146_3_R0_clk),
    .R0_data(mem_146_3_R0_data),
    .R0_en(mem_146_3_R0_en),
    .W0_addr(mem_146_3_W0_addr),
    .W0_clk(mem_146_3_W0_clk),
    .W0_data(mem_146_3_W0_data),
    .W0_en(mem_146_3_W0_en),
    .W0_mask(mem_146_3_W0_mask)
  );
  split_mem_0_ext mem_146_4 (
    .R0_addr(mem_146_4_R0_addr),
    .R0_clk(mem_146_4_R0_clk),
    .R0_data(mem_146_4_R0_data),
    .R0_en(mem_146_4_R0_en),
    .W0_addr(mem_146_4_W0_addr),
    .W0_clk(mem_146_4_W0_clk),
    .W0_data(mem_146_4_W0_data),
    .W0_en(mem_146_4_W0_en),
    .W0_mask(mem_146_4_W0_mask)
  );
  split_mem_0_ext mem_146_5 (
    .R0_addr(mem_146_5_R0_addr),
    .R0_clk(mem_146_5_R0_clk),
    .R0_data(mem_146_5_R0_data),
    .R0_en(mem_146_5_R0_en),
    .W0_addr(mem_146_5_W0_addr),
    .W0_clk(mem_146_5_W0_clk),
    .W0_data(mem_146_5_W0_data),
    .W0_en(mem_146_5_W0_en),
    .W0_mask(mem_146_5_W0_mask)
  );
  split_mem_0_ext mem_146_6 (
    .R0_addr(mem_146_6_R0_addr),
    .R0_clk(mem_146_6_R0_clk),
    .R0_data(mem_146_6_R0_data),
    .R0_en(mem_146_6_R0_en),
    .W0_addr(mem_146_6_W0_addr),
    .W0_clk(mem_146_6_W0_clk),
    .W0_data(mem_146_6_W0_data),
    .W0_en(mem_146_6_W0_en),
    .W0_mask(mem_146_6_W0_mask)
  );
  split_mem_0_ext mem_146_7 (
    .R0_addr(mem_146_7_R0_addr),
    .R0_clk(mem_146_7_R0_clk),
    .R0_data(mem_146_7_R0_data),
    .R0_en(mem_146_7_R0_en),
    .W0_addr(mem_146_7_W0_addr),
    .W0_clk(mem_146_7_W0_clk),
    .W0_data(mem_146_7_W0_data),
    .W0_en(mem_146_7_W0_en),
    .W0_mask(mem_146_7_W0_mask)
  );
  split_mem_0_ext mem_147_0 (
    .R0_addr(mem_147_0_R0_addr),
    .R0_clk(mem_147_0_R0_clk),
    .R0_data(mem_147_0_R0_data),
    .R0_en(mem_147_0_R0_en),
    .W0_addr(mem_147_0_W0_addr),
    .W0_clk(mem_147_0_W0_clk),
    .W0_data(mem_147_0_W0_data),
    .W0_en(mem_147_0_W0_en),
    .W0_mask(mem_147_0_W0_mask)
  );
  split_mem_0_ext mem_147_1 (
    .R0_addr(mem_147_1_R0_addr),
    .R0_clk(mem_147_1_R0_clk),
    .R0_data(mem_147_1_R0_data),
    .R0_en(mem_147_1_R0_en),
    .W0_addr(mem_147_1_W0_addr),
    .W0_clk(mem_147_1_W0_clk),
    .W0_data(mem_147_1_W0_data),
    .W0_en(mem_147_1_W0_en),
    .W0_mask(mem_147_1_W0_mask)
  );
  split_mem_0_ext mem_147_2 (
    .R0_addr(mem_147_2_R0_addr),
    .R0_clk(mem_147_2_R0_clk),
    .R0_data(mem_147_2_R0_data),
    .R0_en(mem_147_2_R0_en),
    .W0_addr(mem_147_2_W0_addr),
    .W0_clk(mem_147_2_W0_clk),
    .W0_data(mem_147_2_W0_data),
    .W0_en(mem_147_2_W0_en),
    .W0_mask(mem_147_2_W0_mask)
  );
  split_mem_0_ext mem_147_3 (
    .R0_addr(mem_147_3_R0_addr),
    .R0_clk(mem_147_3_R0_clk),
    .R0_data(mem_147_3_R0_data),
    .R0_en(mem_147_3_R0_en),
    .W0_addr(mem_147_3_W0_addr),
    .W0_clk(mem_147_3_W0_clk),
    .W0_data(mem_147_3_W0_data),
    .W0_en(mem_147_3_W0_en),
    .W0_mask(mem_147_3_W0_mask)
  );
  split_mem_0_ext mem_147_4 (
    .R0_addr(mem_147_4_R0_addr),
    .R0_clk(mem_147_4_R0_clk),
    .R0_data(mem_147_4_R0_data),
    .R0_en(mem_147_4_R0_en),
    .W0_addr(mem_147_4_W0_addr),
    .W0_clk(mem_147_4_W0_clk),
    .W0_data(mem_147_4_W0_data),
    .W0_en(mem_147_4_W0_en),
    .W0_mask(mem_147_4_W0_mask)
  );
  split_mem_0_ext mem_147_5 (
    .R0_addr(mem_147_5_R0_addr),
    .R0_clk(mem_147_5_R0_clk),
    .R0_data(mem_147_5_R0_data),
    .R0_en(mem_147_5_R0_en),
    .W0_addr(mem_147_5_W0_addr),
    .W0_clk(mem_147_5_W0_clk),
    .W0_data(mem_147_5_W0_data),
    .W0_en(mem_147_5_W0_en),
    .W0_mask(mem_147_5_W0_mask)
  );
  split_mem_0_ext mem_147_6 (
    .R0_addr(mem_147_6_R0_addr),
    .R0_clk(mem_147_6_R0_clk),
    .R0_data(mem_147_6_R0_data),
    .R0_en(mem_147_6_R0_en),
    .W0_addr(mem_147_6_W0_addr),
    .W0_clk(mem_147_6_W0_clk),
    .W0_data(mem_147_6_W0_data),
    .W0_en(mem_147_6_W0_en),
    .W0_mask(mem_147_6_W0_mask)
  );
  split_mem_0_ext mem_147_7 (
    .R0_addr(mem_147_7_R0_addr),
    .R0_clk(mem_147_7_R0_clk),
    .R0_data(mem_147_7_R0_data),
    .R0_en(mem_147_7_R0_en),
    .W0_addr(mem_147_7_W0_addr),
    .W0_clk(mem_147_7_W0_clk),
    .W0_data(mem_147_7_W0_data),
    .W0_en(mem_147_7_W0_en),
    .W0_mask(mem_147_7_W0_mask)
  );
  split_mem_0_ext mem_148_0 (
    .R0_addr(mem_148_0_R0_addr),
    .R0_clk(mem_148_0_R0_clk),
    .R0_data(mem_148_0_R0_data),
    .R0_en(mem_148_0_R0_en),
    .W0_addr(mem_148_0_W0_addr),
    .W0_clk(mem_148_0_W0_clk),
    .W0_data(mem_148_0_W0_data),
    .W0_en(mem_148_0_W0_en),
    .W0_mask(mem_148_0_W0_mask)
  );
  split_mem_0_ext mem_148_1 (
    .R0_addr(mem_148_1_R0_addr),
    .R0_clk(mem_148_1_R0_clk),
    .R0_data(mem_148_1_R0_data),
    .R0_en(mem_148_1_R0_en),
    .W0_addr(mem_148_1_W0_addr),
    .W0_clk(mem_148_1_W0_clk),
    .W0_data(mem_148_1_W0_data),
    .W0_en(mem_148_1_W0_en),
    .W0_mask(mem_148_1_W0_mask)
  );
  split_mem_0_ext mem_148_2 (
    .R0_addr(mem_148_2_R0_addr),
    .R0_clk(mem_148_2_R0_clk),
    .R0_data(mem_148_2_R0_data),
    .R0_en(mem_148_2_R0_en),
    .W0_addr(mem_148_2_W0_addr),
    .W0_clk(mem_148_2_W0_clk),
    .W0_data(mem_148_2_W0_data),
    .W0_en(mem_148_2_W0_en),
    .W0_mask(mem_148_2_W0_mask)
  );
  split_mem_0_ext mem_148_3 (
    .R0_addr(mem_148_3_R0_addr),
    .R0_clk(mem_148_3_R0_clk),
    .R0_data(mem_148_3_R0_data),
    .R0_en(mem_148_3_R0_en),
    .W0_addr(mem_148_3_W0_addr),
    .W0_clk(mem_148_3_W0_clk),
    .W0_data(mem_148_3_W0_data),
    .W0_en(mem_148_3_W0_en),
    .W0_mask(mem_148_3_W0_mask)
  );
  split_mem_0_ext mem_148_4 (
    .R0_addr(mem_148_4_R0_addr),
    .R0_clk(mem_148_4_R0_clk),
    .R0_data(mem_148_4_R0_data),
    .R0_en(mem_148_4_R0_en),
    .W0_addr(mem_148_4_W0_addr),
    .W0_clk(mem_148_4_W0_clk),
    .W0_data(mem_148_4_W0_data),
    .W0_en(mem_148_4_W0_en),
    .W0_mask(mem_148_4_W0_mask)
  );
  split_mem_0_ext mem_148_5 (
    .R0_addr(mem_148_5_R0_addr),
    .R0_clk(mem_148_5_R0_clk),
    .R0_data(mem_148_5_R0_data),
    .R0_en(mem_148_5_R0_en),
    .W0_addr(mem_148_5_W0_addr),
    .W0_clk(mem_148_5_W0_clk),
    .W0_data(mem_148_5_W0_data),
    .W0_en(mem_148_5_W0_en),
    .W0_mask(mem_148_5_W0_mask)
  );
  split_mem_0_ext mem_148_6 (
    .R0_addr(mem_148_6_R0_addr),
    .R0_clk(mem_148_6_R0_clk),
    .R0_data(mem_148_6_R0_data),
    .R0_en(mem_148_6_R0_en),
    .W0_addr(mem_148_6_W0_addr),
    .W0_clk(mem_148_6_W0_clk),
    .W0_data(mem_148_6_W0_data),
    .W0_en(mem_148_6_W0_en),
    .W0_mask(mem_148_6_W0_mask)
  );
  split_mem_0_ext mem_148_7 (
    .R0_addr(mem_148_7_R0_addr),
    .R0_clk(mem_148_7_R0_clk),
    .R0_data(mem_148_7_R0_data),
    .R0_en(mem_148_7_R0_en),
    .W0_addr(mem_148_7_W0_addr),
    .W0_clk(mem_148_7_W0_clk),
    .W0_data(mem_148_7_W0_data),
    .W0_en(mem_148_7_W0_en),
    .W0_mask(mem_148_7_W0_mask)
  );
  split_mem_0_ext mem_149_0 (
    .R0_addr(mem_149_0_R0_addr),
    .R0_clk(mem_149_0_R0_clk),
    .R0_data(mem_149_0_R0_data),
    .R0_en(mem_149_0_R0_en),
    .W0_addr(mem_149_0_W0_addr),
    .W0_clk(mem_149_0_W0_clk),
    .W0_data(mem_149_0_W0_data),
    .W0_en(mem_149_0_W0_en),
    .W0_mask(mem_149_0_W0_mask)
  );
  split_mem_0_ext mem_149_1 (
    .R0_addr(mem_149_1_R0_addr),
    .R0_clk(mem_149_1_R0_clk),
    .R0_data(mem_149_1_R0_data),
    .R0_en(mem_149_1_R0_en),
    .W0_addr(mem_149_1_W0_addr),
    .W0_clk(mem_149_1_W0_clk),
    .W0_data(mem_149_1_W0_data),
    .W0_en(mem_149_1_W0_en),
    .W0_mask(mem_149_1_W0_mask)
  );
  split_mem_0_ext mem_149_2 (
    .R0_addr(mem_149_2_R0_addr),
    .R0_clk(mem_149_2_R0_clk),
    .R0_data(mem_149_2_R0_data),
    .R0_en(mem_149_2_R0_en),
    .W0_addr(mem_149_2_W0_addr),
    .W0_clk(mem_149_2_W0_clk),
    .W0_data(mem_149_2_W0_data),
    .W0_en(mem_149_2_W0_en),
    .W0_mask(mem_149_2_W0_mask)
  );
  split_mem_0_ext mem_149_3 (
    .R0_addr(mem_149_3_R0_addr),
    .R0_clk(mem_149_3_R0_clk),
    .R0_data(mem_149_3_R0_data),
    .R0_en(mem_149_3_R0_en),
    .W0_addr(mem_149_3_W0_addr),
    .W0_clk(mem_149_3_W0_clk),
    .W0_data(mem_149_3_W0_data),
    .W0_en(mem_149_3_W0_en),
    .W0_mask(mem_149_3_W0_mask)
  );
  split_mem_0_ext mem_149_4 (
    .R0_addr(mem_149_4_R0_addr),
    .R0_clk(mem_149_4_R0_clk),
    .R0_data(mem_149_4_R0_data),
    .R0_en(mem_149_4_R0_en),
    .W0_addr(mem_149_4_W0_addr),
    .W0_clk(mem_149_4_W0_clk),
    .W0_data(mem_149_4_W0_data),
    .W0_en(mem_149_4_W0_en),
    .W0_mask(mem_149_4_W0_mask)
  );
  split_mem_0_ext mem_149_5 (
    .R0_addr(mem_149_5_R0_addr),
    .R0_clk(mem_149_5_R0_clk),
    .R0_data(mem_149_5_R0_data),
    .R0_en(mem_149_5_R0_en),
    .W0_addr(mem_149_5_W0_addr),
    .W0_clk(mem_149_5_W0_clk),
    .W0_data(mem_149_5_W0_data),
    .W0_en(mem_149_5_W0_en),
    .W0_mask(mem_149_5_W0_mask)
  );
  split_mem_0_ext mem_149_6 (
    .R0_addr(mem_149_6_R0_addr),
    .R0_clk(mem_149_6_R0_clk),
    .R0_data(mem_149_6_R0_data),
    .R0_en(mem_149_6_R0_en),
    .W0_addr(mem_149_6_W0_addr),
    .W0_clk(mem_149_6_W0_clk),
    .W0_data(mem_149_6_W0_data),
    .W0_en(mem_149_6_W0_en),
    .W0_mask(mem_149_6_W0_mask)
  );
  split_mem_0_ext mem_149_7 (
    .R0_addr(mem_149_7_R0_addr),
    .R0_clk(mem_149_7_R0_clk),
    .R0_data(mem_149_7_R0_data),
    .R0_en(mem_149_7_R0_en),
    .W0_addr(mem_149_7_W0_addr),
    .W0_clk(mem_149_7_W0_clk),
    .W0_data(mem_149_7_W0_data),
    .W0_en(mem_149_7_W0_en),
    .W0_mask(mem_149_7_W0_mask)
  );
  split_mem_0_ext mem_150_0 (
    .R0_addr(mem_150_0_R0_addr),
    .R0_clk(mem_150_0_R0_clk),
    .R0_data(mem_150_0_R0_data),
    .R0_en(mem_150_0_R0_en),
    .W0_addr(mem_150_0_W0_addr),
    .W0_clk(mem_150_0_W0_clk),
    .W0_data(mem_150_0_W0_data),
    .W0_en(mem_150_0_W0_en),
    .W0_mask(mem_150_0_W0_mask)
  );
  split_mem_0_ext mem_150_1 (
    .R0_addr(mem_150_1_R0_addr),
    .R0_clk(mem_150_1_R0_clk),
    .R0_data(mem_150_1_R0_data),
    .R0_en(mem_150_1_R0_en),
    .W0_addr(mem_150_1_W0_addr),
    .W0_clk(mem_150_1_W0_clk),
    .W0_data(mem_150_1_W0_data),
    .W0_en(mem_150_1_W0_en),
    .W0_mask(mem_150_1_W0_mask)
  );
  split_mem_0_ext mem_150_2 (
    .R0_addr(mem_150_2_R0_addr),
    .R0_clk(mem_150_2_R0_clk),
    .R0_data(mem_150_2_R0_data),
    .R0_en(mem_150_2_R0_en),
    .W0_addr(mem_150_2_W0_addr),
    .W0_clk(mem_150_2_W0_clk),
    .W0_data(mem_150_2_W0_data),
    .W0_en(mem_150_2_W0_en),
    .W0_mask(mem_150_2_W0_mask)
  );
  split_mem_0_ext mem_150_3 (
    .R0_addr(mem_150_3_R0_addr),
    .R0_clk(mem_150_3_R0_clk),
    .R0_data(mem_150_3_R0_data),
    .R0_en(mem_150_3_R0_en),
    .W0_addr(mem_150_3_W0_addr),
    .W0_clk(mem_150_3_W0_clk),
    .W0_data(mem_150_3_W0_data),
    .W0_en(mem_150_3_W0_en),
    .W0_mask(mem_150_3_W0_mask)
  );
  split_mem_0_ext mem_150_4 (
    .R0_addr(mem_150_4_R0_addr),
    .R0_clk(mem_150_4_R0_clk),
    .R0_data(mem_150_4_R0_data),
    .R0_en(mem_150_4_R0_en),
    .W0_addr(mem_150_4_W0_addr),
    .W0_clk(mem_150_4_W0_clk),
    .W0_data(mem_150_4_W0_data),
    .W0_en(mem_150_4_W0_en),
    .W0_mask(mem_150_4_W0_mask)
  );
  split_mem_0_ext mem_150_5 (
    .R0_addr(mem_150_5_R0_addr),
    .R0_clk(mem_150_5_R0_clk),
    .R0_data(mem_150_5_R0_data),
    .R0_en(mem_150_5_R0_en),
    .W0_addr(mem_150_5_W0_addr),
    .W0_clk(mem_150_5_W0_clk),
    .W0_data(mem_150_5_W0_data),
    .W0_en(mem_150_5_W0_en),
    .W0_mask(mem_150_5_W0_mask)
  );
  split_mem_0_ext mem_150_6 (
    .R0_addr(mem_150_6_R0_addr),
    .R0_clk(mem_150_6_R0_clk),
    .R0_data(mem_150_6_R0_data),
    .R0_en(mem_150_6_R0_en),
    .W0_addr(mem_150_6_W0_addr),
    .W0_clk(mem_150_6_W0_clk),
    .W0_data(mem_150_6_W0_data),
    .W0_en(mem_150_6_W0_en),
    .W0_mask(mem_150_6_W0_mask)
  );
  split_mem_0_ext mem_150_7 (
    .R0_addr(mem_150_7_R0_addr),
    .R0_clk(mem_150_7_R0_clk),
    .R0_data(mem_150_7_R0_data),
    .R0_en(mem_150_7_R0_en),
    .W0_addr(mem_150_7_W0_addr),
    .W0_clk(mem_150_7_W0_clk),
    .W0_data(mem_150_7_W0_data),
    .W0_en(mem_150_7_W0_en),
    .W0_mask(mem_150_7_W0_mask)
  );
  split_mem_0_ext mem_151_0 (
    .R0_addr(mem_151_0_R0_addr),
    .R0_clk(mem_151_0_R0_clk),
    .R0_data(mem_151_0_R0_data),
    .R0_en(mem_151_0_R0_en),
    .W0_addr(mem_151_0_W0_addr),
    .W0_clk(mem_151_0_W0_clk),
    .W0_data(mem_151_0_W0_data),
    .W0_en(mem_151_0_W0_en),
    .W0_mask(mem_151_0_W0_mask)
  );
  split_mem_0_ext mem_151_1 (
    .R0_addr(mem_151_1_R0_addr),
    .R0_clk(mem_151_1_R0_clk),
    .R0_data(mem_151_1_R0_data),
    .R0_en(mem_151_1_R0_en),
    .W0_addr(mem_151_1_W0_addr),
    .W0_clk(mem_151_1_W0_clk),
    .W0_data(mem_151_1_W0_data),
    .W0_en(mem_151_1_W0_en),
    .W0_mask(mem_151_1_W0_mask)
  );
  split_mem_0_ext mem_151_2 (
    .R0_addr(mem_151_2_R0_addr),
    .R0_clk(mem_151_2_R0_clk),
    .R0_data(mem_151_2_R0_data),
    .R0_en(mem_151_2_R0_en),
    .W0_addr(mem_151_2_W0_addr),
    .W0_clk(mem_151_2_W0_clk),
    .W0_data(mem_151_2_W0_data),
    .W0_en(mem_151_2_W0_en),
    .W0_mask(mem_151_2_W0_mask)
  );
  split_mem_0_ext mem_151_3 (
    .R0_addr(mem_151_3_R0_addr),
    .R0_clk(mem_151_3_R0_clk),
    .R0_data(mem_151_3_R0_data),
    .R0_en(mem_151_3_R0_en),
    .W0_addr(mem_151_3_W0_addr),
    .W0_clk(mem_151_3_W0_clk),
    .W0_data(mem_151_3_W0_data),
    .W0_en(mem_151_3_W0_en),
    .W0_mask(mem_151_3_W0_mask)
  );
  split_mem_0_ext mem_151_4 (
    .R0_addr(mem_151_4_R0_addr),
    .R0_clk(mem_151_4_R0_clk),
    .R0_data(mem_151_4_R0_data),
    .R0_en(mem_151_4_R0_en),
    .W0_addr(mem_151_4_W0_addr),
    .W0_clk(mem_151_4_W0_clk),
    .W0_data(mem_151_4_W0_data),
    .W0_en(mem_151_4_W0_en),
    .W0_mask(mem_151_4_W0_mask)
  );
  split_mem_0_ext mem_151_5 (
    .R0_addr(mem_151_5_R0_addr),
    .R0_clk(mem_151_5_R0_clk),
    .R0_data(mem_151_5_R0_data),
    .R0_en(mem_151_5_R0_en),
    .W0_addr(mem_151_5_W0_addr),
    .W0_clk(mem_151_5_W0_clk),
    .W0_data(mem_151_5_W0_data),
    .W0_en(mem_151_5_W0_en),
    .W0_mask(mem_151_5_W0_mask)
  );
  split_mem_0_ext mem_151_6 (
    .R0_addr(mem_151_6_R0_addr),
    .R0_clk(mem_151_6_R0_clk),
    .R0_data(mem_151_6_R0_data),
    .R0_en(mem_151_6_R0_en),
    .W0_addr(mem_151_6_W0_addr),
    .W0_clk(mem_151_6_W0_clk),
    .W0_data(mem_151_6_W0_data),
    .W0_en(mem_151_6_W0_en),
    .W0_mask(mem_151_6_W0_mask)
  );
  split_mem_0_ext mem_151_7 (
    .R0_addr(mem_151_7_R0_addr),
    .R0_clk(mem_151_7_R0_clk),
    .R0_data(mem_151_7_R0_data),
    .R0_en(mem_151_7_R0_en),
    .W0_addr(mem_151_7_W0_addr),
    .W0_clk(mem_151_7_W0_clk),
    .W0_data(mem_151_7_W0_data),
    .W0_en(mem_151_7_W0_en),
    .W0_mask(mem_151_7_W0_mask)
  );
  split_mem_0_ext mem_152_0 (
    .R0_addr(mem_152_0_R0_addr),
    .R0_clk(mem_152_0_R0_clk),
    .R0_data(mem_152_0_R0_data),
    .R0_en(mem_152_0_R0_en),
    .W0_addr(mem_152_0_W0_addr),
    .W0_clk(mem_152_0_W0_clk),
    .W0_data(mem_152_0_W0_data),
    .W0_en(mem_152_0_W0_en),
    .W0_mask(mem_152_0_W0_mask)
  );
  split_mem_0_ext mem_152_1 (
    .R0_addr(mem_152_1_R0_addr),
    .R0_clk(mem_152_1_R0_clk),
    .R0_data(mem_152_1_R0_data),
    .R0_en(mem_152_1_R0_en),
    .W0_addr(mem_152_1_W0_addr),
    .W0_clk(mem_152_1_W0_clk),
    .W0_data(mem_152_1_W0_data),
    .W0_en(mem_152_1_W0_en),
    .W0_mask(mem_152_1_W0_mask)
  );
  split_mem_0_ext mem_152_2 (
    .R0_addr(mem_152_2_R0_addr),
    .R0_clk(mem_152_2_R0_clk),
    .R0_data(mem_152_2_R0_data),
    .R0_en(mem_152_2_R0_en),
    .W0_addr(mem_152_2_W0_addr),
    .W0_clk(mem_152_2_W0_clk),
    .W0_data(mem_152_2_W0_data),
    .W0_en(mem_152_2_W0_en),
    .W0_mask(mem_152_2_W0_mask)
  );
  split_mem_0_ext mem_152_3 (
    .R0_addr(mem_152_3_R0_addr),
    .R0_clk(mem_152_3_R0_clk),
    .R0_data(mem_152_3_R0_data),
    .R0_en(mem_152_3_R0_en),
    .W0_addr(mem_152_3_W0_addr),
    .W0_clk(mem_152_3_W0_clk),
    .W0_data(mem_152_3_W0_data),
    .W0_en(mem_152_3_W0_en),
    .W0_mask(mem_152_3_W0_mask)
  );
  split_mem_0_ext mem_152_4 (
    .R0_addr(mem_152_4_R0_addr),
    .R0_clk(mem_152_4_R0_clk),
    .R0_data(mem_152_4_R0_data),
    .R0_en(mem_152_4_R0_en),
    .W0_addr(mem_152_4_W0_addr),
    .W0_clk(mem_152_4_W0_clk),
    .W0_data(mem_152_4_W0_data),
    .W0_en(mem_152_4_W0_en),
    .W0_mask(mem_152_4_W0_mask)
  );
  split_mem_0_ext mem_152_5 (
    .R0_addr(mem_152_5_R0_addr),
    .R0_clk(mem_152_5_R0_clk),
    .R0_data(mem_152_5_R0_data),
    .R0_en(mem_152_5_R0_en),
    .W0_addr(mem_152_5_W0_addr),
    .W0_clk(mem_152_5_W0_clk),
    .W0_data(mem_152_5_W0_data),
    .W0_en(mem_152_5_W0_en),
    .W0_mask(mem_152_5_W0_mask)
  );
  split_mem_0_ext mem_152_6 (
    .R0_addr(mem_152_6_R0_addr),
    .R0_clk(mem_152_6_R0_clk),
    .R0_data(mem_152_6_R0_data),
    .R0_en(mem_152_6_R0_en),
    .W0_addr(mem_152_6_W0_addr),
    .W0_clk(mem_152_6_W0_clk),
    .W0_data(mem_152_6_W0_data),
    .W0_en(mem_152_6_W0_en),
    .W0_mask(mem_152_6_W0_mask)
  );
  split_mem_0_ext mem_152_7 (
    .R0_addr(mem_152_7_R0_addr),
    .R0_clk(mem_152_7_R0_clk),
    .R0_data(mem_152_7_R0_data),
    .R0_en(mem_152_7_R0_en),
    .W0_addr(mem_152_7_W0_addr),
    .W0_clk(mem_152_7_W0_clk),
    .W0_data(mem_152_7_W0_data),
    .W0_en(mem_152_7_W0_en),
    .W0_mask(mem_152_7_W0_mask)
  );
  split_mem_0_ext mem_153_0 (
    .R0_addr(mem_153_0_R0_addr),
    .R0_clk(mem_153_0_R0_clk),
    .R0_data(mem_153_0_R0_data),
    .R0_en(mem_153_0_R0_en),
    .W0_addr(mem_153_0_W0_addr),
    .W0_clk(mem_153_0_W0_clk),
    .W0_data(mem_153_0_W0_data),
    .W0_en(mem_153_0_W0_en),
    .W0_mask(mem_153_0_W0_mask)
  );
  split_mem_0_ext mem_153_1 (
    .R0_addr(mem_153_1_R0_addr),
    .R0_clk(mem_153_1_R0_clk),
    .R0_data(mem_153_1_R0_data),
    .R0_en(mem_153_1_R0_en),
    .W0_addr(mem_153_1_W0_addr),
    .W0_clk(mem_153_1_W0_clk),
    .W0_data(mem_153_1_W0_data),
    .W0_en(mem_153_1_W0_en),
    .W0_mask(mem_153_1_W0_mask)
  );
  split_mem_0_ext mem_153_2 (
    .R0_addr(mem_153_2_R0_addr),
    .R0_clk(mem_153_2_R0_clk),
    .R0_data(mem_153_2_R0_data),
    .R0_en(mem_153_2_R0_en),
    .W0_addr(mem_153_2_W0_addr),
    .W0_clk(mem_153_2_W0_clk),
    .W0_data(mem_153_2_W0_data),
    .W0_en(mem_153_2_W0_en),
    .W0_mask(mem_153_2_W0_mask)
  );
  split_mem_0_ext mem_153_3 (
    .R0_addr(mem_153_3_R0_addr),
    .R0_clk(mem_153_3_R0_clk),
    .R0_data(mem_153_3_R0_data),
    .R0_en(mem_153_3_R0_en),
    .W0_addr(mem_153_3_W0_addr),
    .W0_clk(mem_153_3_W0_clk),
    .W0_data(mem_153_3_W0_data),
    .W0_en(mem_153_3_W0_en),
    .W0_mask(mem_153_3_W0_mask)
  );
  split_mem_0_ext mem_153_4 (
    .R0_addr(mem_153_4_R0_addr),
    .R0_clk(mem_153_4_R0_clk),
    .R0_data(mem_153_4_R0_data),
    .R0_en(mem_153_4_R0_en),
    .W0_addr(mem_153_4_W0_addr),
    .W0_clk(mem_153_4_W0_clk),
    .W0_data(mem_153_4_W0_data),
    .W0_en(mem_153_4_W0_en),
    .W0_mask(mem_153_4_W0_mask)
  );
  split_mem_0_ext mem_153_5 (
    .R0_addr(mem_153_5_R0_addr),
    .R0_clk(mem_153_5_R0_clk),
    .R0_data(mem_153_5_R0_data),
    .R0_en(mem_153_5_R0_en),
    .W0_addr(mem_153_5_W0_addr),
    .W0_clk(mem_153_5_W0_clk),
    .W0_data(mem_153_5_W0_data),
    .W0_en(mem_153_5_W0_en),
    .W0_mask(mem_153_5_W0_mask)
  );
  split_mem_0_ext mem_153_6 (
    .R0_addr(mem_153_6_R0_addr),
    .R0_clk(mem_153_6_R0_clk),
    .R0_data(mem_153_6_R0_data),
    .R0_en(mem_153_6_R0_en),
    .W0_addr(mem_153_6_W0_addr),
    .W0_clk(mem_153_6_W0_clk),
    .W0_data(mem_153_6_W0_data),
    .W0_en(mem_153_6_W0_en),
    .W0_mask(mem_153_6_W0_mask)
  );
  split_mem_0_ext mem_153_7 (
    .R0_addr(mem_153_7_R0_addr),
    .R0_clk(mem_153_7_R0_clk),
    .R0_data(mem_153_7_R0_data),
    .R0_en(mem_153_7_R0_en),
    .W0_addr(mem_153_7_W0_addr),
    .W0_clk(mem_153_7_W0_clk),
    .W0_data(mem_153_7_W0_data),
    .W0_en(mem_153_7_W0_en),
    .W0_mask(mem_153_7_W0_mask)
  );
  split_mem_0_ext mem_154_0 (
    .R0_addr(mem_154_0_R0_addr),
    .R0_clk(mem_154_0_R0_clk),
    .R0_data(mem_154_0_R0_data),
    .R0_en(mem_154_0_R0_en),
    .W0_addr(mem_154_0_W0_addr),
    .W0_clk(mem_154_0_W0_clk),
    .W0_data(mem_154_0_W0_data),
    .W0_en(mem_154_0_W0_en),
    .W0_mask(mem_154_0_W0_mask)
  );
  split_mem_0_ext mem_154_1 (
    .R0_addr(mem_154_1_R0_addr),
    .R0_clk(mem_154_1_R0_clk),
    .R0_data(mem_154_1_R0_data),
    .R0_en(mem_154_1_R0_en),
    .W0_addr(mem_154_1_W0_addr),
    .W0_clk(mem_154_1_W0_clk),
    .W0_data(mem_154_1_W0_data),
    .W0_en(mem_154_1_W0_en),
    .W0_mask(mem_154_1_W0_mask)
  );
  split_mem_0_ext mem_154_2 (
    .R0_addr(mem_154_2_R0_addr),
    .R0_clk(mem_154_2_R0_clk),
    .R0_data(mem_154_2_R0_data),
    .R0_en(mem_154_2_R0_en),
    .W0_addr(mem_154_2_W0_addr),
    .W0_clk(mem_154_2_W0_clk),
    .W0_data(mem_154_2_W0_data),
    .W0_en(mem_154_2_W0_en),
    .W0_mask(mem_154_2_W0_mask)
  );
  split_mem_0_ext mem_154_3 (
    .R0_addr(mem_154_3_R0_addr),
    .R0_clk(mem_154_3_R0_clk),
    .R0_data(mem_154_3_R0_data),
    .R0_en(mem_154_3_R0_en),
    .W0_addr(mem_154_3_W0_addr),
    .W0_clk(mem_154_3_W0_clk),
    .W0_data(mem_154_3_W0_data),
    .W0_en(mem_154_3_W0_en),
    .W0_mask(mem_154_3_W0_mask)
  );
  split_mem_0_ext mem_154_4 (
    .R0_addr(mem_154_4_R0_addr),
    .R0_clk(mem_154_4_R0_clk),
    .R0_data(mem_154_4_R0_data),
    .R0_en(mem_154_4_R0_en),
    .W0_addr(mem_154_4_W0_addr),
    .W0_clk(mem_154_4_W0_clk),
    .W0_data(mem_154_4_W0_data),
    .W0_en(mem_154_4_W0_en),
    .W0_mask(mem_154_4_W0_mask)
  );
  split_mem_0_ext mem_154_5 (
    .R0_addr(mem_154_5_R0_addr),
    .R0_clk(mem_154_5_R0_clk),
    .R0_data(mem_154_5_R0_data),
    .R0_en(mem_154_5_R0_en),
    .W0_addr(mem_154_5_W0_addr),
    .W0_clk(mem_154_5_W0_clk),
    .W0_data(mem_154_5_W0_data),
    .W0_en(mem_154_5_W0_en),
    .W0_mask(mem_154_5_W0_mask)
  );
  split_mem_0_ext mem_154_6 (
    .R0_addr(mem_154_6_R0_addr),
    .R0_clk(mem_154_6_R0_clk),
    .R0_data(mem_154_6_R0_data),
    .R0_en(mem_154_6_R0_en),
    .W0_addr(mem_154_6_W0_addr),
    .W0_clk(mem_154_6_W0_clk),
    .W0_data(mem_154_6_W0_data),
    .W0_en(mem_154_6_W0_en),
    .W0_mask(mem_154_6_W0_mask)
  );
  split_mem_0_ext mem_154_7 (
    .R0_addr(mem_154_7_R0_addr),
    .R0_clk(mem_154_7_R0_clk),
    .R0_data(mem_154_7_R0_data),
    .R0_en(mem_154_7_R0_en),
    .W0_addr(mem_154_7_W0_addr),
    .W0_clk(mem_154_7_W0_clk),
    .W0_data(mem_154_7_W0_data),
    .W0_en(mem_154_7_W0_en),
    .W0_mask(mem_154_7_W0_mask)
  );
  split_mem_0_ext mem_155_0 (
    .R0_addr(mem_155_0_R0_addr),
    .R0_clk(mem_155_0_R0_clk),
    .R0_data(mem_155_0_R0_data),
    .R0_en(mem_155_0_R0_en),
    .W0_addr(mem_155_0_W0_addr),
    .W0_clk(mem_155_0_W0_clk),
    .W0_data(mem_155_0_W0_data),
    .W0_en(mem_155_0_W0_en),
    .W0_mask(mem_155_0_W0_mask)
  );
  split_mem_0_ext mem_155_1 (
    .R0_addr(mem_155_1_R0_addr),
    .R0_clk(mem_155_1_R0_clk),
    .R0_data(mem_155_1_R0_data),
    .R0_en(mem_155_1_R0_en),
    .W0_addr(mem_155_1_W0_addr),
    .W0_clk(mem_155_1_W0_clk),
    .W0_data(mem_155_1_W0_data),
    .W0_en(mem_155_1_W0_en),
    .W0_mask(mem_155_1_W0_mask)
  );
  split_mem_0_ext mem_155_2 (
    .R0_addr(mem_155_2_R0_addr),
    .R0_clk(mem_155_2_R0_clk),
    .R0_data(mem_155_2_R0_data),
    .R0_en(mem_155_2_R0_en),
    .W0_addr(mem_155_2_W0_addr),
    .W0_clk(mem_155_2_W0_clk),
    .W0_data(mem_155_2_W0_data),
    .W0_en(mem_155_2_W0_en),
    .W0_mask(mem_155_2_W0_mask)
  );
  split_mem_0_ext mem_155_3 (
    .R0_addr(mem_155_3_R0_addr),
    .R0_clk(mem_155_3_R0_clk),
    .R0_data(mem_155_3_R0_data),
    .R0_en(mem_155_3_R0_en),
    .W0_addr(mem_155_3_W0_addr),
    .W0_clk(mem_155_3_W0_clk),
    .W0_data(mem_155_3_W0_data),
    .W0_en(mem_155_3_W0_en),
    .W0_mask(mem_155_3_W0_mask)
  );
  split_mem_0_ext mem_155_4 (
    .R0_addr(mem_155_4_R0_addr),
    .R0_clk(mem_155_4_R0_clk),
    .R0_data(mem_155_4_R0_data),
    .R0_en(mem_155_4_R0_en),
    .W0_addr(mem_155_4_W0_addr),
    .W0_clk(mem_155_4_W0_clk),
    .W0_data(mem_155_4_W0_data),
    .W0_en(mem_155_4_W0_en),
    .W0_mask(mem_155_4_W0_mask)
  );
  split_mem_0_ext mem_155_5 (
    .R0_addr(mem_155_5_R0_addr),
    .R0_clk(mem_155_5_R0_clk),
    .R0_data(mem_155_5_R0_data),
    .R0_en(mem_155_5_R0_en),
    .W0_addr(mem_155_5_W0_addr),
    .W0_clk(mem_155_5_W0_clk),
    .W0_data(mem_155_5_W0_data),
    .W0_en(mem_155_5_W0_en),
    .W0_mask(mem_155_5_W0_mask)
  );
  split_mem_0_ext mem_155_6 (
    .R0_addr(mem_155_6_R0_addr),
    .R0_clk(mem_155_6_R0_clk),
    .R0_data(mem_155_6_R0_data),
    .R0_en(mem_155_6_R0_en),
    .W0_addr(mem_155_6_W0_addr),
    .W0_clk(mem_155_6_W0_clk),
    .W0_data(mem_155_6_W0_data),
    .W0_en(mem_155_6_W0_en),
    .W0_mask(mem_155_6_W0_mask)
  );
  split_mem_0_ext mem_155_7 (
    .R0_addr(mem_155_7_R0_addr),
    .R0_clk(mem_155_7_R0_clk),
    .R0_data(mem_155_7_R0_data),
    .R0_en(mem_155_7_R0_en),
    .W0_addr(mem_155_7_W0_addr),
    .W0_clk(mem_155_7_W0_clk),
    .W0_data(mem_155_7_W0_data),
    .W0_en(mem_155_7_W0_en),
    .W0_mask(mem_155_7_W0_mask)
  );
  split_mem_0_ext mem_156_0 (
    .R0_addr(mem_156_0_R0_addr),
    .R0_clk(mem_156_0_R0_clk),
    .R0_data(mem_156_0_R0_data),
    .R0_en(mem_156_0_R0_en),
    .W0_addr(mem_156_0_W0_addr),
    .W0_clk(mem_156_0_W0_clk),
    .W0_data(mem_156_0_W0_data),
    .W0_en(mem_156_0_W0_en),
    .W0_mask(mem_156_0_W0_mask)
  );
  split_mem_0_ext mem_156_1 (
    .R0_addr(mem_156_1_R0_addr),
    .R0_clk(mem_156_1_R0_clk),
    .R0_data(mem_156_1_R0_data),
    .R0_en(mem_156_1_R0_en),
    .W0_addr(mem_156_1_W0_addr),
    .W0_clk(mem_156_1_W0_clk),
    .W0_data(mem_156_1_W0_data),
    .W0_en(mem_156_1_W0_en),
    .W0_mask(mem_156_1_W0_mask)
  );
  split_mem_0_ext mem_156_2 (
    .R0_addr(mem_156_2_R0_addr),
    .R0_clk(mem_156_2_R0_clk),
    .R0_data(mem_156_2_R0_data),
    .R0_en(mem_156_2_R0_en),
    .W0_addr(mem_156_2_W0_addr),
    .W0_clk(mem_156_2_W0_clk),
    .W0_data(mem_156_2_W0_data),
    .W0_en(mem_156_2_W0_en),
    .W0_mask(mem_156_2_W0_mask)
  );
  split_mem_0_ext mem_156_3 (
    .R0_addr(mem_156_3_R0_addr),
    .R0_clk(mem_156_3_R0_clk),
    .R0_data(mem_156_3_R0_data),
    .R0_en(mem_156_3_R0_en),
    .W0_addr(mem_156_3_W0_addr),
    .W0_clk(mem_156_3_W0_clk),
    .W0_data(mem_156_3_W0_data),
    .W0_en(mem_156_3_W0_en),
    .W0_mask(mem_156_3_W0_mask)
  );
  split_mem_0_ext mem_156_4 (
    .R0_addr(mem_156_4_R0_addr),
    .R0_clk(mem_156_4_R0_clk),
    .R0_data(mem_156_4_R0_data),
    .R0_en(mem_156_4_R0_en),
    .W0_addr(mem_156_4_W0_addr),
    .W0_clk(mem_156_4_W0_clk),
    .W0_data(mem_156_4_W0_data),
    .W0_en(mem_156_4_W0_en),
    .W0_mask(mem_156_4_W0_mask)
  );
  split_mem_0_ext mem_156_5 (
    .R0_addr(mem_156_5_R0_addr),
    .R0_clk(mem_156_5_R0_clk),
    .R0_data(mem_156_5_R0_data),
    .R0_en(mem_156_5_R0_en),
    .W0_addr(mem_156_5_W0_addr),
    .W0_clk(mem_156_5_W0_clk),
    .W0_data(mem_156_5_W0_data),
    .W0_en(mem_156_5_W0_en),
    .W0_mask(mem_156_5_W0_mask)
  );
  split_mem_0_ext mem_156_6 (
    .R0_addr(mem_156_6_R0_addr),
    .R0_clk(mem_156_6_R0_clk),
    .R0_data(mem_156_6_R0_data),
    .R0_en(mem_156_6_R0_en),
    .W0_addr(mem_156_6_W0_addr),
    .W0_clk(mem_156_6_W0_clk),
    .W0_data(mem_156_6_W0_data),
    .W0_en(mem_156_6_W0_en),
    .W0_mask(mem_156_6_W0_mask)
  );
  split_mem_0_ext mem_156_7 (
    .R0_addr(mem_156_7_R0_addr),
    .R0_clk(mem_156_7_R0_clk),
    .R0_data(mem_156_7_R0_data),
    .R0_en(mem_156_7_R0_en),
    .W0_addr(mem_156_7_W0_addr),
    .W0_clk(mem_156_7_W0_clk),
    .W0_data(mem_156_7_W0_data),
    .W0_en(mem_156_7_W0_en),
    .W0_mask(mem_156_7_W0_mask)
  );
  split_mem_0_ext mem_157_0 (
    .R0_addr(mem_157_0_R0_addr),
    .R0_clk(mem_157_0_R0_clk),
    .R0_data(mem_157_0_R0_data),
    .R0_en(mem_157_0_R0_en),
    .W0_addr(mem_157_0_W0_addr),
    .W0_clk(mem_157_0_W0_clk),
    .W0_data(mem_157_0_W0_data),
    .W0_en(mem_157_0_W0_en),
    .W0_mask(mem_157_0_W0_mask)
  );
  split_mem_0_ext mem_157_1 (
    .R0_addr(mem_157_1_R0_addr),
    .R0_clk(mem_157_1_R0_clk),
    .R0_data(mem_157_1_R0_data),
    .R0_en(mem_157_1_R0_en),
    .W0_addr(mem_157_1_W0_addr),
    .W0_clk(mem_157_1_W0_clk),
    .W0_data(mem_157_1_W0_data),
    .W0_en(mem_157_1_W0_en),
    .W0_mask(mem_157_1_W0_mask)
  );
  split_mem_0_ext mem_157_2 (
    .R0_addr(mem_157_2_R0_addr),
    .R0_clk(mem_157_2_R0_clk),
    .R0_data(mem_157_2_R0_data),
    .R0_en(mem_157_2_R0_en),
    .W0_addr(mem_157_2_W0_addr),
    .W0_clk(mem_157_2_W0_clk),
    .W0_data(mem_157_2_W0_data),
    .W0_en(mem_157_2_W0_en),
    .W0_mask(mem_157_2_W0_mask)
  );
  split_mem_0_ext mem_157_3 (
    .R0_addr(mem_157_3_R0_addr),
    .R0_clk(mem_157_3_R0_clk),
    .R0_data(mem_157_3_R0_data),
    .R0_en(mem_157_3_R0_en),
    .W0_addr(mem_157_3_W0_addr),
    .W0_clk(mem_157_3_W0_clk),
    .W0_data(mem_157_3_W0_data),
    .W0_en(mem_157_3_W0_en),
    .W0_mask(mem_157_3_W0_mask)
  );
  split_mem_0_ext mem_157_4 (
    .R0_addr(mem_157_4_R0_addr),
    .R0_clk(mem_157_4_R0_clk),
    .R0_data(mem_157_4_R0_data),
    .R0_en(mem_157_4_R0_en),
    .W0_addr(mem_157_4_W0_addr),
    .W0_clk(mem_157_4_W0_clk),
    .W0_data(mem_157_4_W0_data),
    .W0_en(mem_157_4_W0_en),
    .W0_mask(mem_157_4_W0_mask)
  );
  split_mem_0_ext mem_157_5 (
    .R0_addr(mem_157_5_R0_addr),
    .R0_clk(mem_157_5_R0_clk),
    .R0_data(mem_157_5_R0_data),
    .R0_en(mem_157_5_R0_en),
    .W0_addr(mem_157_5_W0_addr),
    .W0_clk(mem_157_5_W0_clk),
    .W0_data(mem_157_5_W0_data),
    .W0_en(mem_157_5_W0_en),
    .W0_mask(mem_157_5_W0_mask)
  );
  split_mem_0_ext mem_157_6 (
    .R0_addr(mem_157_6_R0_addr),
    .R0_clk(mem_157_6_R0_clk),
    .R0_data(mem_157_6_R0_data),
    .R0_en(mem_157_6_R0_en),
    .W0_addr(mem_157_6_W0_addr),
    .W0_clk(mem_157_6_W0_clk),
    .W0_data(mem_157_6_W0_data),
    .W0_en(mem_157_6_W0_en),
    .W0_mask(mem_157_6_W0_mask)
  );
  split_mem_0_ext mem_157_7 (
    .R0_addr(mem_157_7_R0_addr),
    .R0_clk(mem_157_7_R0_clk),
    .R0_data(mem_157_7_R0_data),
    .R0_en(mem_157_7_R0_en),
    .W0_addr(mem_157_7_W0_addr),
    .W0_clk(mem_157_7_W0_clk),
    .W0_data(mem_157_7_W0_data),
    .W0_en(mem_157_7_W0_en),
    .W0_mask(mem_157_7_W0_mask)
  );
  split_mem_0_ext mem_158_0 (
    .R0_addr(mem_158_0_R0_addr),
    .R0_clk(mem_158_0_R0_clk),
    .R0_data(mem_158_0_R0_data),
    .R0_en(mem_158_0_R0_en),
    .W0_addr(mem_158_0_W0_addr),
    .W0_clk(mem_158_0_W0_clk),
    .W0_data(mem_158_0_W0_data),
    .W0_en(mem_158_0_W0_en),
    .W0_mask(mem_158_0_W0_mask)
  );
  split_mem_0_ext mem_158_1 (
    .R0_addr(mem_158_1_R0_addr),
    .R0_clk(mem_158_1_R0_clk),
    .R0_data(mem_158_1_R0_data),
    .R0_en(mem_158_1_R0_en),
    .W0_addr(mem_158_1_W0_addr),
    .W0_clk(mem_158_1_W0_clk),
    .W0_data(mem_158_1_W0_data),
    .W0_en(mem_158_1_W0_en),
    .W0_mask(mem_158_1_W0_mask)
  );
  split_mem_0_ext mem_158_2 (
    .R0_addr(mem_158_2_R0_addr),
    .R0_clk(mem_158_2_R0_clk),
    .R0_data(mem_158_2_R0_data),
    .R0_en(mem_158_2_R0_en),
    .W0_addr(mem_158_2_W0_addr),
    .W0_clk(mem_158_2_W0_clk),
    .W0_data(mem_158_2_W0_data),
    .W0_en(mem_158_2_W0_en),
    .W0_mask(mem_158_2_W0_mask)
  );
  split_mem_0_ext mem_158_3 (
    .R0_addr(mem_158_3_R0_addr),
    .R0_clk(mem_158_3_R0_clk),
    .R0_data(mem_158_3_R0_data),
    .R0_en(mem_158_3_R0_en),
    .W0_addr(mem_158_3_W0_addr),
    .W0_clk(mem_158_3_W0_clk),
    .W0_data(mem_158_3_W0_data),
    .W0_en(mem_158_3_W0_en),
    .W0_mask(mem_158_3_W0_mask)
  );
  split_mem_0_ext mem_158_4 (
    .R0_addr(mem_158_4_R0_addr),
    .R0_clk(mem_158_4_R0_clk),
    .R0_data(mem_158_4_R0_data),
    .R0_en(mem_158_4_R0_en),
    .W0_addr(mem_158_4_W0_addr),
    .W0_clk(mem_158_4_W0_clk),
    .W0_data(mem_158_4_W0_data),
    .W0_en(mem_158_4_W0_en),
    .W0_mask(mem_158_4_W0_mask)
  );
  split_mem_0_ext mem_158_5 (
    .R0_addr(mem_158_5_R0_addr),
    .R0_clk(mem_158_5_R0_clk),
    .R0_data(mem_158_5_R0_data),
    .R0_en(mem_158_5_R0_en),
    .W0_addr(mem_158_5_W0_addr),
    .W0_clk(mem_158_5_W0_clk),
    .W0_data(mem_158_5_W0_data),
    .W0_en(mem_158_5_W0_en),
    .W0_mask(mem_158_5_W0_mask)
  );
  split_mem_0_ext mem_158_6 (
    .R0_addr(mem_158_6_R0_addr),
    .R0_clk(mem_158_6_R0_clk),
    .R0_data(mem_158_6_R0_data),
    .R0_en(mem_158_6_R0_en),
    .W0_addr(mem_158_6_W0_addr),
    .W0_clk(mem_158_6_W0_clk),
    .W0_data(mem_158_6_W0_data),
    .W0_en(mem_158_6_W0_en),
    .W0_mask(mem_158_6_W0_mask)
  );
  split_mem_0_ext mem_158_7 (
    .R0_addr(mem_158_7_R0_addr),
    .R0_clk(mem_158_7_R0_clk),
    .R0_data(mem_158_7_R0_data),
    .R0_en(mem_158_7_R0_en),
    .W0_addr(mem_158_7_W0_addr),
    .W0_clk(mem_158_7_W0_clk),
    .W0_data(mem_158_7_W0_data),
    .W0_en(mem_158_7_W0_en),
    .W0_mask(mem_158_7_W0_mask)
  );
  split_mem_0_ext mem_159_0 (
    .R0_addr(mem_159_0_R0_addr),
    .R0_clk(mem_159_0_R0_clk),
    .R0_data(mem_159_0_R0_data),
    .R0_en(mem_159_0_R0_en),
    .W0_addr(mem_159_0_W0_addr),
    .W0_clk(mem_159_0_W0_clk),
    .W0_data(mem_159_0_W0_data),
    .W0_en(mem_159_0_W0_en),
    .W0_mask(mem_159_0_W0_mask)
  );
  split_mem_0_ext mem_159_1 (
    .R0_addr(mem_159_1_R0_addr),
    .R0_clk(mem_159_1_R0_clk),
    .R0_data(mem_159_1_R0_data),
    .R0_en(mem_159_1_R0_en),
    .W0_addr(mem_159_1_W0_addr),
    .W0_clk(mem_159_1_W0_clk),
    .W0_data(mem_159_1_W0_data),
    .W0_en(mem_159_1_W0_en),
    .W0_mask(mem_159_1_W0_mask)
  );
  split_mem_0_ext mem_159_2 (
    .R0_addr(mem_159_2_R0_addr),
    .R0_clk(mem_159_2_R0_clk),
    .R0_data(mem_159_2_R0_data),
    .R0_en(mem_159_2_R0_en),
    .W0_addr(mem_159_2_W0_addr),
    .W0_clk(mem_159_2_W0_clk),
    .W0_data(mem_159_2_W0_data),
    .W0_en(mem_159_2_W0_en),
    .W0_mask(mem_159_2_W0_mask)
  );
  split_mem_0_ext mem_159_3 (
    .R0_addr(mem_159_3_R0_addr),
    .R0_clk(mem_159_3_R0_clk),
    .R0_data(mem_159_3_R0_data),
    .R0_en(mem_159_3_R0_en),
    .W0_addr(mem_159_3_W0_addr),
    .W0_clk(mem_159_3_W0_clk),
    .W0_data(mem_159_3_W0_data),
    .W0_en(mem_159_3_W0_en),
    .W0_mask(mem_159_3_W0_mask)
  );
  split_mem_0_ext mem_159_4 (
    .R0_addr(mem_159_4_R0_addr),
    .R0_clk(mem_159_4_R0_clk),
    .R0_data(mem_159_4_R0_data),
    .R0_en(mem_159_4_R0_en),
    .W0_addr(mem_159_4_W0_addr),
    .W0_clk(mem_159_4_W0_clk),
    .W0_data(mem_159_4_W0_data),
    .W0_en(mem_159_4_W0_en),
    .W0_mask(mem_159_4_W0_mask)
  );
  split_mem_0_ext mem_159_5 (
    .R0_addr(mem_159_5_R0_addr),
    .R0_clk(mem_159_5_R0_clk),
    .R0_data(mem_159_5_R0_data),
    .R0_en(mem_159_5_R0_en),
    .W0_addr(mem_159_5_W0_addr),
    .W0_clk(mem_159_5_W0_clk),
    .W0_data(mem_159_5_W0_data),
    .W0_en(mem_159_5_W0_en),
    .W0_mask(mem_159_5_W0_mask)
  );
  split_mem_0_ext mem_159_6 (
    .R0_addr(mem_159_6_R0_addr),
    .R0_clk(mem_159_6_R0_clk),
    .R0_data(mem_159_6_R0_data),
    .R0_en(mem_159_6_R0_en),
    .W0_addr(mem_159_6_W0_addr),
    .W0_clk(mem_159_6_W0_clk),
    .W0_data(mem_159_6_W0_data),
    .W0_en(mem_159_6_W0_en),
    .W0_mask(mem_159_6_W0_mask)
  );
  split_mem_0_ext mem_159_7 (
    .R0_addr(mem_159_7_R0_addr),
    .R0_clk(mem_159_7_R0_clk),
    .R0_data(mem_159_7_R0_data),
    .R0_en(mem_159_7_R0_en),
    .W0_addr(mem_159_7_W0_addr),
    .W0_clk(mem_159_7_W0_clk),
    .W0_data(mem_159_7_W0_data),
    .W0_en(mem_159_7_W0_en),
    .W0_mask(mem_159_7_W0_mask)
  );
  split_mem_0_ext mem_160_0 (
    .R0_addr(mem_160_0_R0_addr),
    .R0_clk(mem_160_0_R0_clk),
    .R0_data(mem_160_0_R0_data),
    .R0_en(mem_160_0_R0_en),
    .W0_addr(mem_160_0_W0_addr),
    .W0_clk(mem_160_0_W0_clk),
    .W0_data(mem_160_0_W0_data),
    .W0_en(mem_160_0_W0_en),
    .W0_mask(mem_160_0_W0_mask)
  );
  split_mem_0_ext mem_160_1 (
    .R0_addr(mem_160_1_R0_addr),
    .R0_clk(mem_160_1_R0_clk),
    .R0_data(mem_160_1_R0_data),
    .R0_en(mem_160_1_R0_en),
    .W0_addr(mem_160_1_W0_addr),
    .W0_clk(mem_160_1_W0_clk),
    .W0_data(mem_160_1_W0_data),
    .W0_en(mem_160_1_W0_en),
    .W0_mask(mem_160_1_W0_mask)
  );
  split_mem_0_ext mem_160_2 (
    .R0_addr(mem_160_2_R0_addr),
    .R0_clk(mem_160_2_R0_clk),
    .R0_data(mem_160_2_R0_data),
    .R0_en(mem_160_2_R0_en),
    .W0_addr(mem_160_2_W0_addr),
    .W0_clk(mem_160_2_W0_clk),
    .W0_data(mem_160_2_W0_data),
    .W0_en(mem_160_2_W0_en),
    .W0_mask(mem_160_2_W0_mask)
  );
  split_mem_0_ext mem_160_3 (
    .R0_addr(mem_160_3_R0_addr),
    .R0_clk(mem_160_3_R0_clk),
    .R0_data(mem_160_3_R0_data),
    .R0_en(mem_160_3_R0_en),
    .W0_addr(mem_160_3_W0_addr),
    .W0_clk(mem_160_3_W0_clk),
    .W0_data(mem_160_3_W0_data),
    .W0_en(mem_160_3_W0_en),
    .W0_mask(mem_160_3_W0_mask)
  );
  split_mem_0_ext mem_160_4 (
    .R0_addr(mem_160_4_R0_addr),
    .R0_clk(mem_160_4_R0_clk),
    .R0_data(mem_160_4_R0_data),
    .R0_en(mem_160_4_R0_en),
    .W0_addr(mem_160_4_W0_addr),
    .W0_clk(mem_160_4_W0_clk),
    .W0_data(mem_160_4_W0_data),
    .W0_en(mem_160_4_W0_en),
    .W0_mask(mem_160_4_W0_mask)
  );
  split_mem_0_ext mem_160_5 (
    .R0_addr(mem_160_5_R0_addr),
    .R0_clk(mem_160_5_R0_clk),
    .R0_data(mem_160_5_R0_data),
    .R0_en(mem_160_5_R0_en),
    .W0_addr(mem_160_5_W0_addr),
    .W0_clk(mem_160_5_W0_clk),
    .W0_data(mem_160_5_W0_data),
    .W0_en(mem_160_5_W0_en),
    .W0_mask(mem_160_5_W0_mask)
  );
  split_mem_0_ext mem_160_6 (
    .R0_addr(mem_160_6_R0_addr),
    .R0_clk(mem_160_6_R0_clk),
    .R0_data(mem_160_6_R0_data),
    .R0_en(mem_160_6_R0_en),
    .W0_addr(mem_160_6_W0_addr),
    .W0_clk(mem_160_6_W0_clk),
    .W0_data(mem_160_6_W0_data),
    .W0_en(mem_160_6_W0_en),
    .W0_mask(mem_160_6_W0_mask)
  );
  split_mem_0_ext mem_160_7 (
    .R0_addr(mem_160_7_R0_addr),
    .R0_clk(mem_160_7_R0_clk),
    .R0_data(mem_160_7_R0_data),
    .R0_en(mem_160_7_R0_en),
    .W0_addr(mem_160_7_W0_addr),
    .W0_clk(mem_160_7_W0_clk),
    .W0_data(mem_160_7_W0_data),
    .W0_en(mem_160_7_W0_en),
    .W0_mask(mem_160_7_W0_mask)
  );
  split_mem_0_ext mem_161_0 (
    .R0_addr(mem_161_0_R0_addr),
    .R0_clk(mem_161_0_R0_clk),
    .R0_data(mem_161_0_R0_data),
    .R0_en(mem_161_0_R0_en),
    .W0_addr(mem_161_0_W0_addr),
    .W0_clk(mem_161_0_W0_clk),
    .W0_data(mem_161_0_W0_data),
    .W0_en(mem_161_0_W0_en),
    .W0_mask(mem_161_0_W0_mask)
  );
  split_mem_0_ext mem_161_1 (
    .R0_addr(mem_161_1_R0_addr),
    .R0_clk(mem_161_1_R0_clk),
    .R0_data(mem_161_1_R0_data),
    .R0_en(mem_161_1_R0_en),
    .W0_addr(mem_161_1_W0_addr),
    .W0_clk(mem_161_1_W0_clk),
    .W0_data(mem_161_1_W0_data),
    .W0_en(mem_161_1_W0_en),
    .W0_mask(mem_161_1_W0_mask)
  );
  split_mem_0_ext mem_161_2 (
    .R0_addr(mem_161_2_R0_addr),
    .R0_clk(mem_161_2_R0_clk),
    .R0_data(mem_161_2_R0_data),
    .R0_en(mem_161_2_R0_en),
    .W0_addr(mem_161_2_W0_addr),
    .W0_clk(mem_161_2_W0_clk),
    .W0_data(mem_161_2_W0_data),
    .W0_en(mem_161_2_W0_en),
    .W0_mask(mem_161_2_W0_mask)
  );
  split_mem_0_ext mem_161_3 (
    .R0_addr(mem_161_3_R0_addr),
    .R0_clk(mem_161_3_R0_clk),
    .R0_data(mem_161_3_R0_data),
    .R0_en(mem_161_3_R0_en),
    .W0_addr(mem_161_3_W0_addr),
    .W0_clk(mem_161_3_W0_clk),
    .W0_data(mem_161_3_W0_data),
    .W0_en(mem_161_3_W0_en),
    .W0_mask(mem_161_3_W0_mask)
  );
  split_mem_0_ext mem_161_4 (
    .R0_addr(mem_161_4_R0_addr),
    .R0_clk(mem_161_4_R0_clk),
    .R0_data(mem_161_4_R0_data),
    .R0_en(mem_161_4_R0_en),
    .W0_addr(mem_161_4_W0_addr),
    .W0_clk(mem_161_4_W0_clk),
    .W0_data(mem_161_4_W0_data),
    .W0_en(mem_161_4_W0_en),
    .W0_mask(mem_161_4_W0_mask)
  );
  split_mem_0_ext mem_161_5 (
    .R0_addr(mem_161_5_R0_addr),
    .R0_clk(mem_161_5_R0_clk),
    .R0_data(mem_161_5_R0_data),
    .R0_en(mem_161_5_R0_en),
    .W0_addr(mem_161_5_W0_addr),
    .W0_clk(mem_161_5_W0_clk),
    .W0_data(mem_161_5_W0_data),
    .W0_en(mem_161_5_W0_en),
    .W0_mask(mem_161_5_W0_mask)
  );
  split_mem_0_ext mem_161_6 (
    .R0_addr(mem_161_6_R0_addr),
    .R0_clk(mem_161_6_R0_clk),
    .R0_data(mem_161_6_R0_data),
    .R0_en(mem_161_6_R0_en),
    .W0_addr(mem_161_6_W0_addr),
    .W0_clk(mem_161_6_W0_clk),
    .W0_data(mem_161_6_W0_data),
    .W0_en(mem_161_6_W0_en),
    .W0_mask(mem_161_6_W0_mask)
  );
  split_mem_0_ext mem_161_7 (
    .R0_addr(mem_161_7_R0_addr),
    .R0_clk(mem_161_7_R0_clk),
    .R0_data(mem_161_7_R0_data),
    .R0_en(mem_161_7_R0_en),
    .W0_addr(mem_161_7_W0_addr),
    .W0_clk(mem_161_7_W0_clk),
    .W0_data(mem_161_7_W0_data),
    .W0_en(mem_161_7_W0_en),
    .W0_mask(mem_161_7_W0_mask)
  );
  split_mem_0_ext mem_162_0 (
    .R0_addr(mem_162_0_R0_addr),
    .R0_clk(mem_162_0_R0_clk),
    .R0_data(mem_162_0_R0_data),
    .R0_en(mem_162_0_R0_en),
    .W0_addr(mem_162_0_W0_addr),
    .W0_clk(mem_162_0_W0_clk),
    .W0_data(mem_162_0_W0_data),
    .W0_en(mem_162_0_W0_en),
    .W0_mask(mem_162_0_W0_mask)
  );
  split_mem_0_ext mem_162_1 (
    .R0_addr(mem_162_1_R0_addr),
    .R0_clk(mem_162_1_R0_clk),
    .R0_data(mem_162_1_R0_data),
    .R0_en(mem_162_1_R0_en),
    .W0_addr(mem_162_1_W0_addr),
    .W0_clk(mem_162_1_W0_clk),
    .W0_data(mem_162_1_W0_data),
    .W0_en(mem_162_1_W0_en),
    .W0_mask(mem_162_1_W0_mask)
  );
  split_mem_0_ext mem_162_2 (
    .R0_addr(mem_162_2_R0_addr),
    .R0_clk(mem_162_2_R0_clk),
    .R0_data(mem_162_2_R0_data),
    .R0_en(mem_162_2_R0_en),
    .W0_addr(mem_162_2_W0_addr),
    .W0_clk(mem_162_2_W0_clk),
    .W0_data(mem_162_2_W0_data),
    .W0_en(mem_162_2_W0_en),
    .W0_mask(mem_162_2_W0_mask)
  );
  split_mem_0_ext mem_162_3 (
    .R0_addr(mem_162_3_R0_addr),
    .R0_clk(mem_162_3_R0_clk),
    .R0_data(mem_162_3_R0_data),
    .R0_en(mem_162_3_R0_en),
    .W0_addr(mem_162_3_W0_addr),
    .W0_clk(mem_162_3_W0_clk),
    .W0_data(mem_162_3_W0_data),
    .W0_en(mem_162_3_W0_en),
    .W0_mask(mem_162_3_W0_mask)
  );
  split_mem_0_ext mem_162_4 (
    .R0_addr(mem_162_4_R0_addr),
    .R0_clk(mem_162_4_R0_clk),
    .R0_data(mem_162_4_R0_data),
    .R0_en(mem_162_4_R0_en),
    .W0_addr(mem_162_4_W0_addr),
    .W0_clk(mem_162_4_W0_clk),
    .W0_data(mem_162_4_W0_data),
    .W0_en(mem_162_4_W0_en),
    .W0_mask(mem_162_4_W0_mask)
  );
  split_mem_0_ext mem_162_5 (
    .R0_addr(mem_162_5_R0_addr),
    .R0_clk(mem_162_5_R0_clk),
    .R0_data(mem_162_5_R0_data),
    .R0_en(mem_162_5_R0_en),
    .W0_addr(mem_162_5_W0_addr),
    .W0_clk(mem_162_5_W0_clk),
    .W0_data(mem_162_5_W0_data),
    .W0_en(mem_162_5_W0_en),
    .W0_mask(mem_162_5_W0_mask)
  );
  split_mem_0_ext mem_162_6 (
    .R0_addr(mem_162_6_R0_addr),
    .R0_clk(mem_162_6_R0_clk),
    .R0_data(mem_162_6_R0_data),
    .R0_en(mem_162_6_R0_en),
    .W0_addr(mem_162_6_W0_addr),
    .W0_clk(mem_162_6_W0_clk),
    .W0_data(mem_162_6_W0_data),
    .W0_en(mem_162_6_W0_en),
    .W0_mask(mem_162_6_W0_mask)
  );
  split_mem_0_ext mem_162_7 (
    .R0_addr(mem_162_7_R0_addr),
    .R0_clk(mem_162_7_R0_clk),
    .R0_data(mem_162_7_R0_data),
    .R0_en(mem_162_7_R0_en),
    .W0_addr(mem_162_7_W0_addr),
    .W0_clk(mem_162_7_W0_clk),
    .W0_data(mem_162_7_W0_data),
    .W0_en(mem_162_7_W0_en),
    .W0_mask(mem_162_7_W0_mask)
  );
  split_mem_0_ext mem_163_0 (
    .R0_addr(mem_163_0_R0_addr),
    .R0_clk(mem_163_0_R0_clk),
    .R0_data(mem_163_0_R0_data),
    .R0_en(mem_163_0_R0_en),
    .W0_addr(mem_163_0_W0_addr),
    .W0_clk(mem_163_0_W0_clk),
    .W0_data(mem_163_0_W0_data),
    .W0_en(mem_163_0_W0_en),
    .W0_mask(mem_163_0_W0_mask)
  );
  split_mem_0_ext mem_163_1 (
    .R0_addr(mem_163_1_R0_addr),
    .R0_clk(mem_163_1_R0_clk),
    .R0_data(mem_163_1_R0_data),
    .R0_en(mem_163_1_R0_en),
    .W0_addr(mem_163_1_W0_addr),
    .W0_clk(mem_163_1_W0_clk),
    .W0_data(mem_163_1_W0_data),
    .W0_en(mem_163_1_W0_en),
    .W0_mask(mem_163_1_W0_mask)
  );
  split_mem_0_ext mem_163_2 (
    .R0_addr(mem_163_2_R0_addr),
    .R0_clk(mem_163_2_R0_clk),
    .R0_data(mem_163_2_R0_data),
    .R0_en(mem_163_2_R0_en),
    .W0_addr(mem_163_2_W0_addr),
    .W0_clk(mem_163_2_W0_clk),
    .W0_data(mem_163_2_W0_data),
    .W0_en(mem_163_2_W0_en),
    .W0_mask(mem_163_2_W0_mask)
  );
  split_mem_0_ext mem_163_3 (
    .R0_addr(mem_163_3_R0_addr),
    .R0_clk(mem_163_3_R0_clk),
    .R0_data(mem_163_3_R0_data),
    .R0_en(mem_163_3_R0_en),
    .W0_addr(mem_163_3_W0_addr),
    .W0_clk(mem_163_3_W0_clk),
    .W0_data(mem_163_3_W0_data),
    .W0_en(mem_163_3_W0_en),
    .W0_mask(mem_163_3_W0_mask)
  );
  split_mem_0_ext mem_163_4 (
    .R0_addr(mem_163_4_R0_addr),
    .R0_clk(mem_163_4_R0_clk),
    .R0_data(mem_163_4_R0_data),
    .R0_en(mem_163_4_R0_en),
    .W0_addr(mem_163_4_W0_addr),
    .W0_clk(mem_163_4_W0_clk),
    .W0_data(mem_163_4_W0_data),
    .W0_en(mem_163_4_W0_en),
    .W0_mask(mem_163_4_W0_mask)
  );
  split_mem_0_ext mem_163_5 (
    .R0_addr(mem_163_5_R0_addr),
    .R0_clk(mem_163_5_R0_clk),
    .R0_data(mem_163_5_R0_data),
    .R0_en(mem_163_5_R0_en),
    .W0_addr(mem_163_5_W0_addr),
    .W0_clk(mem_163_5_W0_clk),
    .W0_data(mem_163_5_W0_data),
    .W0_en(mem_163_5_W0_en),
    .W0_mask(mem_163_5_W0_mask)
  );
  split_mem_0_ext mem_163_6 (
    .R0_addr(mem_163_6_R0_addr),
    .R0_clk(mem_163_6_R0_clk),
    .R0_data(mem_163_6_R0_data),
    .R0_en(mem_163_6_R0_en),
    .W0_addr(mem_163_6_W0_addr),
    .W0_clk(mem_163_6_W0_clk),
    .W0_data(mem_163_6_W0_data),
    .W0_en(mem_163_6_W0_en),
    .W0_mask(mem_163_6_W0_mask)
  );
  split_mem_0_ext mem_163_7 (
    .R0_addr(mem_163_7_R0_addr),
    .R0_clk(mem_163_7_R0_clk),
    .R0_data(mem_163_7_R0_data),
    .R0_en(mem_163_7_R0_en),
    .W0_addr(mem_163_7_W0_addr),
    .W0_clk(mem_163_7_W0_clk),
    .W0_data(mem_163_7_W0_data),
    .W0_en(mem_163_7_W0_en),
    .W0_mask(mem_163_7_W0_mask)
  );
  split_mem_0_ext mem_164_0 (
    .R0_addr(mem_164_0_R0_addr),
    .R0_clk(mem_164_0_R0_clk),
    .R0_data(mem_164_0_R0_data),
    .R0_en(mem_164_0_R0_en),
    .W0_addr(mem_164_0_W0_addr),
    .W0_clk(mem_164_0_W0_clk),
    .W0_data(mem_164_0_W0_data),
    .W0_en(mem_164_0_W0_en),
    .W0_mask(mem_164_0_W0_mask)
  );
  split_mem_0_ext mem_164_1 (
    .R0_addr(mem_164_1_R0_addr),
    .R0_clk(mem_164_1_R0_clk),
    .R0_data(mem_164_1_R0_data),
    .R0_en(mem_164_1_R0_en),
    .W0_addr(mem_164_1_W0_addr),
    .W0_clk(mem_164_1_W0_clk),
    .W0_data(mem_164_1_W0_data),
    .W0_en(mem_164_1_W0_en),
    .W0_mask(mem_164_1_W0_mask)
  );
  split_mem_0_ext mem_164_2 (
    .R0_addr(mem_164_2_R0_addr),
    .R0_clk(mem_164_2_R0_clk),
    .R0_data(mem_164_2_R0_data),
    .R0_en(mem_164_2_R0_en),
    .W0_addr(mem_164_2_W0_addr),
    .W0_clk(mem_164_2_W0_clk),
    .W0_data(mem_164_2_W0_data),
    .W0_en(mem_164_2_W0_en),
    .W0_mask(mem_164_2_W0_mask)
  );
  split_mem_0_ext mem_164_3 (
    .R0_addr(mem_164_3_R0_addr),
    .R0_clk(mem_164_3_R0_clk),
    .R0_data(mem_164_3_R0_data),
    .R0_en(mem_164_3_R0_en),
    .W0_addr(mem_164_3_W0_addr),
    .W0_clk(mem_164_3_W0_clk),
    .W0_data(mem_164_3_W0_data),
    .W0_en(mem_164_3_W0_en),
    .W0_mask(mem_164_3_W0_mask)
  );
  split_mem_0_ext mem_164_4 (
    .R0_addr(mem_164_4_R0_addr),
    .R0_clk(mem_164_4_R0_clk),
    .R0_data(mem_164_4_R0_data),
    .R0_en(mem_164_4_R0_en),
    .W0_addr(mem_164_4_W0_addr),
    .W0_clk(mem_164_4_W0_clk),
    .W0_data(mem_164_4_W0_data),
    .W0_en(mem_164_4_W0_en),
    .W0_mask(mem_164_4_W0_mask)
  );
  split_mem_0_ext mem_164_5 (
    .R0_addr(mem_164_5_R0_addr),
    .R0_clk(mem_164_5_R0_clk),
    .R0_data(mem_164_5_R0_data),
    .R0_en(mem_164_5_R0_en),
    .W0_addr(mem_164_5_W0_addr),
    .W0_clk(mem_164_5_W0_clk),
    .W0_data(mem_164_5_W0_data),
    .W0_en(mem_164_5_W0_en),
    .W0_mask(mem_164_5_W0_mask)
  );
  split_mem_0_ext mem_164_6 (
    .R0_addr(mem_164_6_R0_addr),
    .R0_clk(mem_164_6_R0_clk),
    .R0_data(mem_164_6_R0_data),
    .R0_en(mem_164_6_R0_en),
    .W0_addr(mem_164_6_W0_addr),
    .W0_clk(mem_164_6_W0_clk),
    .W0_data(mem_164_6_W0_data),
    .W0_en(mem_164_6_W0_en),
    .W0_mask(mem_164_6_W0_mask)
  );
  split_mem_0_ext mem_164_7 (
    .R0_addr(mem_164_7_R0_addr),
    .R0_clk(mem_164_7_R0_clk),
    .R0_data(mem_164_7_R0_data),
    .R0_en(mem_164_7_R0_en),
    .W0_addr(mem_164_7_W0_addr),
    .W0_clk(mem_164_7_W0_clk),
    .W0_data(mem_164_7_W0_data),
    .W0_en(mem_164_7_W0_en),
    .W0_mask(mem_164_7_W0_mask)
  );
  split_mem_0_ext mem_165_0 (
    .R0_addr(mem_165_0_R0_addr),
    .R0_clk(mem_165_0_R0_clk),
    .R0_data(mem_165_0_R0_data),
    .R0_en(mem_165_0_R0_en),
    .W0_addr(mem_165_0_W0_addr),
    .W0_clk(mem_165_0_W0_clk),
    .W0_data(mem_165_0_W0_data),
    .W0_en(mem_165_0_W0_en),
    .W0_mask(mem_165_0_W0_mask)
  );
  split_mem_0_ext mem_165_1 (
    .R0_addr(mem_165_1_R0_addr),
    .R0_clk(mem_165_1_R0_clk),
    .R0_data(mem_165_1_R0_data),
    .R0_en(mem_165_1_R0_en),
    .W0_addr(mem_165_1_W0_addr),
    .W0_clk(mem_165_1_W0_clk),
    .W0_data(mem_165_1_W0_data),
    .W0_en(mem_165_1_W0_en),
    .W0_mask(mem_165_1_W0_mask)
  );
  split_mem_0_ext mem_165_2 (
    .R0_addr(mem_165_2_R0_addr),
    .R0_clk(mem_165_2_R0_clk),
    .R0_data(mem_165_2_R0_data),
    .R0_en(mem_165_2_R0_en),
    .W0_addr(mem_165_2_W0_addr),
    .W0_clk(mem_165_2_W0_clk),
    .W0_data(mem_165_2_W0_data),
    .W0_en(mem_165_2_W0_en),
    .W0_mask(mem_165_2_W0_mask)
  );
  split_mem_0_ext mem_165_3 (
    .R0_addr(mem_165_3_R0_addr),
    .R0_clk(mem_165_3_R0_clk),
    .R0_data(mem_165_3_R0_data),
    .R0_en(mem_165_3_R0_en),
    .W0_addr(mem_165_3_W0_addr),
    .W0_clk(mem_165_3_W0_clk),
    .W0_data(mem_165_3_W0_data),
    .W0_en(mem_165_3_W0_en),
    .W0_mask(mem_165_3_W0_mask)
  );
  split_mem_0_ext mem_165_4 (
    .R0_addr(mem_165_4_R0_addr),
    .R0_clk(mem_165_4_R0_clk),
    .R0_data(mem_165_4_R0_data),
    .R0_en(mem_165_4_R0_en),
    .W0_addr(mem_165_4_W0_addr),
    .W0_clk(mem_165_4_W0_clk),
    .W0_data(mem_165_4_W0_data),
    .W0_en(mem_165_4_W0_en),
    .W0_mask(mem_165_4_W0_mask)
  );
  split_mem_0_ext mem_165_5 (
    .R0_addr(mem_165_5_R0_addr),
    .R0_clk(mem_165_5_R0_clk),
    .R0_data(mem_165_5_R0_data),
    .R0_en(mem_165_5_R0_en),
    .W0_addr(mem_165_5_W0_addr),
    .W0_clk(mem_165_5_W0_clk),
    .W0_data(mem_165_5_W0_data),
    .W0_en(mem_165_5_W0_en),
    .W0_mask(mem_165_5_W0_mask)
  );
  split_mem_0_ext mem_165_6 (
    .R0_addr(mem_165_6_R0_addr),
    .R0_clk(mem_165_6_R0_clk),
    .R0_data(mem_165_6_R0_data),
    .R0_en(mem_165_6_R0_en),
    .W0_addr(mem_165_6_W0_addr),
    .W0_clk(mem_165_6_W0_clk),
    .W0_data(mem_165_6_W0_data),
    .W0_en(mem_165_6_W0_en),
    .W0_mask(mem_165_6_W0_mask)
  );
  split_mem_0_ext mem_165_7 (
    .R0_addr(mem_165_7_R0_addr),
    .R0_clk(mem_165_7_R0_clk),
    .R0_data(mem_165_7_R0_data),
    .R0_en(mem_165_7_R0_en),
    .W0_addr(mem_165_7_W0_addr),
    .W0_clk(mem_165_7_W0_clk),
    .W0_data(mem_165_7_W0_data),
    .W0_en(mem_165_7_W0_en),
    .W0_mask(mem_165_7_W0_mask)
  );
  split_mem_0_ext mem_166_0 (
    .R0_addr(mem_166_0_R0_addr),
    .R0_clk(mem_166_0_R0_clk),
    .R0_data(mem_166_0_R0_data),
    .R0_en(mem_166_0_R0_en),
    .W0_addr(mem_166_0_W0_addr),
    .W0_clk(mem_166_0_W0_clk),
    .W0_data(mem_166_0_W0_data),
    .W0_en(mem_166_0_W0_en),
    .W0_mask(mem_166_0_W0_mask)
  );
  split_mem_0_ext mem_166_1 (
    .R0_addr(mem_166_1_R0_addr),
    .R0_clk(mem_166_1_R0_clk),
    .R0_data(mem_166_1_R0_data),
    .R0_en(mem_166_1_R0_en),
    .W0_addr(mem_166_1_W0_addr),
    .W0_clk(mem_166_1_W0_clk),
    .W0_data(mem_166_1_W0_data),
    .W0_en(mem_166_1_W0_en),
    .W0_mask(mem_166_1_W0_mask)
  );
  split_mem_0_ext mem_166_2 (
    .R0_addr(mem_166_2_R0_addr),
    .R0_clk(mem_166_2_R0_clk),
    .R0_data(mem_166_2_R0_data),
    .R0_en(mem_166_2_R0_en),
    .W0_addr(mem_166_2_W0_addr),
    .W0_clk(mem_166_2_W0_clk),
    .W0_data(mem_166_2_W0_data),
    .W0_en(mem_166_2_W0_en),
    .W0_mask(mem_166_2_W0_mask)
  );
  split_mem_0_ext mem_166_3 (
    .R0_addr(mem_166_3_R0_addr),
    .R0_clk(mem_166_3_R0_clk),
    .R0_data(mem_166_3_R0_data),
    .R0_en(mem_166_3_R0_en),
    .W0_addr(mem_166_3_W0_addr),
    .W0_clk(mem_166_3_W0_clk),
    .W0_data(mem_166_3_W0_data),
    .W0_en(mem_166_3_W0_en),
    .W0_mask(mem_166_3_W0_mask)
  );
  split_mem_0_ext mem_166_4 (
    .R0_addr(mem_166_4_R0_addr),
    .R0_clk(mem_166_4_R0_clk),
    .R0_data(mem_166_4_R0_data),
    .R0_en(mem_166_4_R0_en),
    .W0_addr(mem_166_4_W0_addr),
    .W0_clk(mem_166_4_W0_clk),
    .W0_data(mem_166_4_W0_data),
    .W0_en(mem_166_4_W0_en),
    .W0_mask(mem_166_4_W0_mask)
  );
  split_mem_0_ext mem_166_5 (
    .R0_addr(mem_166_5_R0_addr),
    .R0_clk(mem_166_5_R0_clk),
    .R0_data(mem_166_5_R0_data),
    .R0_en(mem_166_5_R0_en),
    .W0_addr(mem_166_5_W0_addr),
    .W0_clk(mem_166_5_W0_clk),
    .W0_data(mem_166_5_W0_data),
    .W0_en(mem_166_5_W0_en),
    .W0_mask(mem_166_5_W0_mask)
  );
  split_mem_0_ext mem_166_6 (
    .R0_addr(mem_166_6_R0_addr),
    .R0_clk(mem_166_6_R0_clk),
    .R0_data(mem_166_6_R0_data),
    .R0_en(mem_166_6_R0_en),
    .W0_addr(mem_166_6_W0_addr),
    .W0_clk(mem_166_6_W0_clk),
    .W0_data(mem_166_6_W0_data),
    .W0_en(mem_166_6_W0_en),
    .W0_mask(mem_166_6_W0_mask)
  );
  split_mem_0_ext mem_166_7 (
    .R0_addr(mem_166_7_R0_addr),
    .R0_clk(mem_166_7_R0_clk),
    .R0_data(mem_166_7_R0_data),
    .R0_en(mem_166_7_R0_en),
    .W0_addr(mem_166_7_W0_addr),
    .W0_clk(mem_166_7_W0_clk),
    .W0_data(mem_166_7_W0_data),
    .W0_en(mem_166_7_W0_en),
    .W0_mask(mem_166_7_W0_mask)
  );
  split_mem_0_ext mem_167_0 (
    .R0_addr(mem_167_0_R0_addr),
    .R0_clk(mem_167_0_R0_clk),
    .R0_data(mem_167_0_R0_data),
    .R0_en(mem_167_0_R0_en),
    .W0_addr(mem_167_0_W0_addr),
    .W0_clk(mem_167_0_W0_clk),
    .W0_data(mem_167_0_W0_data),
    .W0_en(mem_167_0_W0_en),
    .W0_mask(mem_167_0_W0_mask)
  );
  split_mem_0_ext mem_167_1 (
    .R0_addr(mem_167_1_R0_addr),
    .R0_clk(mem_167_1_R0_clk),
    .R0_data(mem_167_1_R0_data),
    .R0_en(mem_167_1_R0_en),
    .W0_addr(mem_167_1_W0_addr),
    .W0_clk(mem_167_1_W0_clk),
    .W0_data(mem_167_1_W0_data),
    .W0_en(mem_167_1_W0_en),
    .W0_mask(mem_167_1_W0_mask)
  );
  split_mem_0_ext mem_167_2 (
    .R0_addr(mem_167_2_R0_addr),
    .R0_clk(mem_167_2_R0_clk),
    .R0_data(mem_167_2_R0_data),
    .R0_en(mem_167_2_R0_en),
    .W0_addr(mem_167_2_W0_addr),
    .W0_clk(mem_167_2_W0_clk),
    .W0_data(mem_167_2_W0_data),
    .W0_en(mem_167_2_W0_en),
    .W0_mask(mem_167_2_W0_mask)
  );
  split_mem_0_ext mem_167_3 (
    .R0_addr(mem_167_3_R0_addr),
    .R0_clk(mem_167_3_R0_clk),
    .R0_data(mem_167_3_R0_data),
    .R0_en(mem_167_3_R0_en),
    .W0_addr(mem_167_3_W0_addr),
    .W0_clk(mem_167_3_W0_clk),
    .W0_data(mem_167_3_W0_data),
    .W0_en(mem_167_3_W0_en),
    .W0_mask(mem_167_3_W0_mask)
  );
  split_mem_0_ext mem_167_4 (
    .R0_addr(mem_167_4_R0_addr),
    .R0_clk(mem_167_4_R0_clk),
    .R0_data(mem_167_4_R0_data),
    .R0_en(mem_167_4_R0_en),
    .W0_addr(mem_167_4_W0_addr),
    .W0_clk(mem_167_4_W0_clk),
    .W0_data(mem_167_4_W0_data),
    .W0_en(mem_167_4_W0_en),
    .W0_mask(mem_167_4_W0_mask)
  );
  split_mem_0_ext mem_167_5 (
    .R0_addr(mem_167_5_R0_addr),
    .R0_clk(mem_167_5_R0_clk),
    .R0_data(mem_167_5_R0_data),
    .R0_en(mem_167_5_R0_en),
    .W0_addr(mem_167_5_W0_addr),
    .W0_clk(mem_167_5_W0_clk),
    .W0_data(mem_167_5_W0_data),
    .W0_en(mem_167_5_W0_en),
    .W0_mask(mem_167_5_W0_mask)
  );
  split_mem_0_ext mem_167_6 (
    .R0_addr(mem_167_6_R0_addr),
    .R0_clk(mem_167_6_R0_clk),
    .R0_data(mem_167_6_R0_data),
    .R0_en(mem_167_6_R0_en),
    .W0_addr(mem_167_6_W0_addr),
    .W0_clk(mem_167_6_W0_clk),
    .W0_data(mem_167_6_W0_data),
    .W0_en(mem_167_6_W0_en),
    .W0_mask(mem_167_6_W0_mask)
  );
  split_mem_0_ext mem_167_7 (
    .R0_addr(mem_167_7_R0_addr),
    .R0_clk(mem_167_7_R0_clk),
    .R0_data(mem_167_7_R0_data),
    .R0_en(mem_167_7_R0_en),
    .W0_addr(mem_167_7_W0_addr),
    .W0_clk(mem_167_7_W0_clk),
    .W0_data(mem_167_7_W0_data),
    .W0_en(mem_167_7_W0_en),
    .W0_mask(mem_167_7_W0_mask)
  );
  split_mem_0_ext mem_168_0 (
    .R0_addr(mem_168_0_R0_addr),
    .R0_clk(mem_168_0_R0_clk),
    .R0_data(mem_168_0_R0_data),
    .R0_en(mem_168_0_R0_en),
    .W0_addr(mem_168_0_W0_addr),
    .W0_clk(mem_168_0_W0_clk),
    .W0_data(mem_168_0_W0_data),
    .W0_en(mem_168_0_W0_en),
    .W0_mask(mem_168_0_W0_mask)
  );
  split_mem_0_ext mem_168_1 (
    .R0_addr(mem_168_1_R0_addr),
    .R0_clk(mem_168_1_R0_clk),
    .R0_data(mem_168_1_R0_data),
    .R0_en(mem_168_1_R0_en),
    .W0_addr(mem_168_1_W0_addr),
    .W0_clk(mem_168_1_W0_clk),
    .W0_data(mem_168_1_W0_data),
    .W0_en(mem_168_1_W0_en),
    .W0_mask(mem_168_1_W0_mask)
  );
  split_mem_0_ext mem_168_2 (
    .R0_addr(mem_168_2_R0_addr),
    .R0_clk(mem_168_2_R0_clk),
    .R0_data(mem_168_2_R0_data),
    .R0_en(mem_168_2_R0_en),
    .W0_addr(mem_168_2_W0_addr),
    .W0_clk(mem_168_2_W0_clk),
    .W0_data(mem_168_2_W0_data),
    .W0_en(mem_168_2_W0_en),
    .W0_mask(mem_168_2_W0_mask)
  );
  split_mem_0_ext mem_168_3 (
    .R0_addr(mem_168_3_R0_addr),
    .R0_clk(mem_168_3_R0_clk),
    .R0_data(mem_168_3_R0_data),
    .R0_en(mem_168_3_R0_en),
    .W0_addr(mem_168_3_W0_addr),
    .W0_clk(mem_168_3_W0_clk),
    .W0_data(mem_168_3_W0_data),
    .W0_en(mem_168_3_W0_en),
    .W0_mask(mem_168_3_W0_mask)
  );
  split_mem_0_ext mem_168_4 (
    .R0_addr(mem_168_4_R0_addr),
    .R0_clk(mem_168_4_R0_clk),
    .R0_data(mem_168_4_R0_data),
    .R0_en(mem_168_4_R0_en),
    .W0_addr(mem_168_4_W0_addr),
    .W0_clk(mem_168_4_W0_clk),
    .W0_data(mem_168_4_W0_data),
    .W0_en(mem_168_4_W0_en),
    .W0_mask(mem_168_4_W0_mask)
  );
  split_mem_0_ext mem_168_5 (
    .R0_addr(mem_168_5_R0_addr),
    .R0_clk(mem_168_5_R0_clk),
    .R0_data(mem_168_5_R0_data),
    .R0_en(mem_168_5_R0_en),
    .W0_addr(mem_168_5_W0_addr),
    .W0_clk(mem_168_5_W0_clk),
    .W0_data(mem_168_5_W0_data),
    .W0_en(mem_168_5_W0_en),
    .W0_mask(mem_168_5_W0_mask)
  );
  split_mem_0_ext mem_168_6 (
    .R0_addr(mem_168_6_R0_addr),
    .R0_clk(mem_168_6_R0_clk),
    .R0_data(mem_168_6_R0_data),
    .R0_en(mem_168_6_R0_en),
    .W0_addr(mem_168_6_W0_addr),
    .W0_clk(mem_168_6_W0_clk),
    .W0_data(mem_168_6_W0_data),
    .W0_en(mem_168_6_W0_en),
    .W0_mask(mem_168_6_W0_mask)
  );
  split_mem_0_ext mem_168_7 (
    .R0_addr(mem_168_7_R0_addr),
    .R0_clk(mem_168_7_R0_clk),
    .R0_data(mem_168_7_R0_data),
    .R0_en(mem_168_7_R0_en),
    .W0_addr(mem_168_7_W0_addr),
    .W0_clk(mem_168_7_W0_clk),
    .W0_data(mem_168_7_W0_data),
    .W0_en(mem_168_7_W0_en),
    .W0_mask(mem_168_7_W0_mask)
  );
  split_mem_0_ext mem_169_0 (
    .R0_addr(mem_169_0_R0_addr),
    .R0_clk(mem_169_0_R0_clk),
    .R0_data(mem_169_0_R0_data),
    .R0_en(mem_169_0_R0_en),
    .W0_addr(mem_169_0_W0_addr),
    .W0_clk(mem_169_0_W0_clk),
    .W0_data(mem_169_0_W0_data),
    .W0_en(mem_169_0_W0_en),
    .W0_mask(mem_169_0_W0_mask)
  );
  split_mem_0_ext mem_169_1 (
    .R0_addr(mem_169_1_R0_addr),
    .R0_clk(mem_169_1_R0_clk),
    .R0_data(mem_169_1_R0_data),
    .R0_en(mem_169_1_R0_en),
    .W0_addr(mem_169_1_W0_addr),
    .W0_clk(mem_169_1_W0_clk),
    .W0_data(mem_169_1_W0_data),
    .W0_en(mem_169_1_W0_en),
    .W0_mask(mem_169_1_W0_mask)
  );
  split_mem_0_ext mem_169_2 (
    .R0_addr(mem_169_2_R0_addr),
    .R0_clk(mem_169_2_R0_clk),
    .R0_data(mem_169_2_R0_data),
    .R0_en(mem_169_2_R0_en),
    .W0_addr(mem_169_2_W0_addr),
    .W0_clk(mem_169_2_W0_clk),
    .W0_data(mem_169_2_W0_data),
    .W0_en(mem_169_2_W0_en),
    .W0_mask(mem_169_2_W0_mask)
  );
  split_mem_0_ext mem_169_3 (
    .R0_addr(mem_169_3_R0_addr),
    .R0_clk(mem_169_3_R0_clk),
    .R0_data(mem_169_3_R0_data),
    .R0_en(mem_169_3_R0_en),
    .W0_addr(mem_169_3_W0_addr),
    .W0_clk(mem_169_3_W0_clk),
    .W0_data(mem_169_3_W0_data),
    .W0_en(mem_169_3_W0_en),
    .W0_mask(mem_169_3_W0_mask)
  );
  split_mem_0_ext mem_169_4 (
    .R0_addr(mem_169_4_R0_addr),
    .R0_clk(mem_169_4_R0_clk),
    .R0_data(mem_169_4_R0_data),
    .R0_en(mem_169_4_R0_en),
    .W0_addr(mem_169_4_W0_addr),
    .W0_clk(mem_169_4_W0_clk),
    .W0_data(mem_169_4_W0_data),
    .W0_en(mem_169_4_W0_en),
    .W0_mask(mem_169_4_W0_mask)
  );
  split_mem_0_ext mem_169_5 (
    .R0_addr(mem_169_5_R0_addr),
    .R0_clk(mem_169_5_R0_clk),
    .R0_data(mem_169_5_R0_data),
    .R0_en(mem_169_5_R0_en),
    .W0_addr(mem_169_5_W0_addr),
    .W0_clk(mem_169_5_W0_clk),
    .W0_data(mem_169_5_W0_data),
    .W0_en(mem_169_5_W0_en),
    .W0_mask(mem_169_5_W0_mask)
  );
  split_mem_0_ext mem_169_6 (
    .R0_addr(mem_169_6_R0_addr),
    .R0_clk(mem_169_6_R0_clk),
    .R0_data(mem_169_6_R0_data),
    .R0_en(mem_169_6_R0_en),
    .W0_addr(mem_169_6_W0_addr),
    .W0_clk(mem_169_6_W0_clk),
    .W0_data(mem_169_6_W0_data),
    .W0_en(mem_169_6_W0_en),
    .W0_mask(mem_169_6_W0_mask)
  );
  split_mem_0_ext mem_169_7 (
    .R0_addr(mem_169_7_R0_addr),
    .R0_clk(mem_169_7_R0_clk),
    .R0_data(mem_169_7_R0_data),
    .R0_en(mem_169_7_R0_en),
    .W0_addr(mem_169_7_W0_addr),
    .W0_clk(mem_169_7_W0_clk),
    .W0_data(mem_169_7_W0_data),
    .W0_en(mem_169_7_W0_en),
    .W0_mask(mem_169_7_W0_mask)
  );
  split_mem_0_ext mem_170_0 (
    .R0_addr(mem_170_0_R0_addr),
    .R0_clk(mem_170_0_R0_clk),
    .R0_data(mem_170_0_R0_data),
    .R0_en(mem_170_0_R0_en),
    .W0_addr(mem_170_0_W0_addr),
    .W0_clk(mem_170_0_W0_clk),
    .W0_data(mem_170_0_W0_data),
    .W0_en(mem_170_0_W0_en),
    .W0_mask(mem_170_0_W0_mask)
  );
  split_mem_0_ext mem_170_1 (
    .R0_addr(mem_170_1_R0_addr),
    .R0_clk(mem_170_1_R0_clk),
    .R0_data(mem_170_1_R0_data),
    .R0_en(mem_170_1_R0_en),
    .W0_addr(mem_170_1_W0_addr),
    .W0_clk(mem_170_1_W0_clk),
    .W0_data(mem_170_1_W0_data),
    .W0_en(mem_170_1_W0_en),
    .W0_mask(mem_170_1_W0_mask)
  );
  split_mem_0_ext mem_170_2 (
    .R0_addr(mem_170_2_R0_addr),
    .R0_clk(mem_170_2_R0_clk),
    .R0_data(mem_170_2_R0_data),
    .R0_en(mem_170_2_R0_en),
    .W0_addr(mem_170_2_W0_addr),
    .W0_clk(mem_170_2_W0_clk),
    .W0_data(mem_170_2_W0_data),
    .W0_en(mem_170_2_W0_en),
    .W0_mask(mem_170_2_W0_mask)
  );
  split_mem_0_ext mem_170_3 (
    .R0_addr(mem_170_3_R0_addr),
    .R0_clk(mem_170_3_R0_clk),
    .R0_data(mem_170_3_R0_data),
    .R0_en(mem_170_3_R0_en),
    .W0_addr(mem_170_3_W0_addr),
    .W0_clk(mem_170_3_W0_clk),
    .W0_data(mem_170_3_W0_data),
    .W0_en(mem_170_3_W0_en),
    .W0_mask(mem_170_3_W0_mask)
  );
  split_mem_0_ext mem_170_4 (
    .R0_addr(mem_170_4_R0_addr),
    .R0_clk(mem_170_4_R0_clk),
    .R0_data(mem_170_4_R0_data),
    .R0_en(mem_170_4_R0_en),
    .W0_addr(mem_170_4_W0_addr),
    .W0_clk(mem_170_4_W0_clk),
    .W0_data(mem_170_4_W0_data),
    .W0_en(mem_170_4_W0_en),
    .W0_mask(mem_170_4_W0_mask)
  );
  split_mem_0_ext mem_170_5 (
    .R0_addr(mem_170_5_R0_addr),
    .R0_clk(mem_170_5_R0_clk),
    .R0_data(mem_170_5_R0_data),
    .R0_en(mem_170_5_R0_en),
    .W0_addr(mem_170_5_W0_addr),
    .W0_clk(mem_170_5_W0_clk),
    .W0_data(mem_170_5_W0_data),
    .W0_en(mem_170_5_W0_en),
    .W0_mask(mem_170_5_W0_mask)
  );
  split_mem_0_ext mem_170_6 (
    .R0_addr(mem_170_6_R0_addr),
    .R0_clk(mem_170_6_R0_clk),
    .R0_data(mem_170_6_R0_data),
    .R0_en(mem_170_6_R0_en),
    .W0_addr(mem_170_6_W0_addr),
    .W0_clk(mem_170_6_W0_clk),
    .W0_data(mem_170_6_W0_data),
    .W0_en(mem_170_6_W0_en),
    .W0_mask(mem_170_6_W0_mask)
  );
  split_mem_0_ext mem_170_7 (
    .R0_addr(mem_170_7_R0_addr),
    .R0_clk(mem_170_7_R0_clk),
    .R0_data(mem_170_7_R0_data),
    .R0_en(mem_170_7_R0_en),
    .W0_addr(mem_170_7_W0_addr),
    .W0_clk(mem_170_7_W0_clk),
    .W0_data(mem_170_7_W0_data),
    .W0_en(mem_170_7_W0_en),
    .W0_mask(mem_170_7_W0_mask)
  );
  split_mem_0_ext mem_171_0 (
    .R0_addr(mem_171_0_R0_addr),
    .R0_clk(mem_171_0_R0_clk),
    .R0_data(mem_171_0_R0_data),
    .R0_en(mem_171_0_R0_en),
    .W0_addr(mem_171_0_W0_addr),
    .W0_clk(mem_171_0_W0_clk),
    .W0_data(mem_171_0_W0_data),
    .W0_en(mem_171_0_W0_en),
    .W0_mask(mem_171_0_W0_mask)
  );
  split_mem_0_ext mem_171_1 (
    .R0_addr(mem_171_1_R0_addr),
    .R0_clk(mem_171_1_R0_clk),
    .R0_data(mem_171_1_R0_data),
    .R0_en(mem_171_1_R0_en),
    .W0_addr(mem_171_1_W0_addr),
    .W0_clk(mem_171_1_W0_clk),
    .W0_data(mem_171_1_W0_data),
    .W0_en(mem_171_1_W0_en),
    .W0_mask(mem_171_1_W0_mask)
  );
  split_mem_0_ext mem_171_2 (
    .R0_addr(mem_171_2_R0_addr),
    .R0_clk(mem_171_2_R0_clk),
    .R0_data(mem_171_2_R0_data),
    .R0_en(mem_171_2_R0_en),
    .W0_addr(mem_171_2_W0_addr),
    .W0_clk(mem_171_2_W0_clk),
    .W0_data(mem_171_2_W0_data),
    .W0_en(mem_171_2_W0_en),
    .W0_mask(mem_171_2_W0_mask)
  );
  split_mem_0_ext mem_171_3 (
    .R0_addr(mem_171_3_R0_addr),
    .R0_clk(mem_171_3_R0_clk),
    .R0_data(mem_171_3_R0_data),
    .R0_en(mem_171_3_R0_en),
    .W0_addr(mem_171_3_W0_addr),
    .W0_clk(mem_171_3_W0_clk),
    .W0_data(mem_171_3_W0_data),
    .W0_en(mem_171_3_W0_en),
    .W0_mask(mem_171_3_W0_mask)
  );
  split_mem_0_ext mem_171_4 (
    .R0_addr(mem_171_4_R0_addr),
    .R0_clk(mem_171_4_R0_clk),
    .R0_data(mem_171_4_R0_data),
    .R0_en(mem_171_4_R0_en),
    .W0_addr(mem_171_4_W0_addr),
    .W0_clk(mem_171_4_W0_clk),
    .W0_data(mem_171_4_W0_data),
    .W0_en(mem_171_4_W0_en),
    .W0_mask(mem_171_4_W0_mask)
  );
  split_mem_0_ext mem_171_5 (
    .R0_addr(mem_171_5_R0_addr),
    .R0_clk(mem_171_5_R0_clk),
    .R0_data(mem_171_5_R0_data),
    .R0_en(mem_171_5_R0_en),
    .W0_addr(mem_171_5_W0_addr),
    .W0_clk(mem_171_5_W0_clk),
    .W0_data(mem_171_5_W0_data),
    .W0_en(mem_171_5_W0_en),
    .W0_mask(mem_171_5_W0_mask)
  );
  split_mem_0_ext mem_171_6 (
    .R0_addr(mem_171_6_R0_addr),
    .R0_clk(mem_171_6_R0_clk),
    .R0_data(mem_171_6_R0_data),
    .R0_en(mem_171_6_R0_en),
    .W0_addr(mem_171_6_W0_addr),
    .W0_clk(mem_171_6_W0_clk),
    .W0_data(mem_171_6_W0_data),
    .W0_en(mem_171_6_W0_en),
    .W0_mask(mem_171_6_W0_mask)
  );
  split_mem_0_ext mem_171_7 (
    .R0_addr(mem_171_7_R0_addr),
    .R0_clk(mem_171_7_R0_clk),
    .R0_data(mem_171_7_R0_data),
    .R0_en(mem_171_7_R0_en),
    .W0_addr(mem_171_7_W0_addr),
    .W0_clk(mem_171_7_W0_clk),
    .W0_data(mem_171_7_W0_data),
    .W0_en(mem_171_7_W0_en),
    .W0_mask(mem_171_7_W0_mask)
  );
  split_mem_0_ext mem_172_0 (
    .R0_addr(mem_172_0_R0_addr),
    .R0_clk(mem_172_0_R0_clk),
    .R0_data(mem_172_0_R0_data),
    .R0_en(mem_172_0_R0_en),
    .W0_addr(mem_172_0_W0_addr),
    .W0_clk(mem_172_0_W0_clk),
    .W0_data(mem_172_0_W0_data),
    .W0_en(mem_172_0_W0_en),
    .W0_mask(mem_172_0_W0_mask)
  );
  split_mem_0_ext mem_172_1 (
    .R0_addr(mem_172_1_R0_addr),
    .R0_clk(mem_172_1_R0_clk),
    .R0_data(mem_172_1_R0_data),
    .R0_en(mem_172_1_R0_en),
    .W0_addr(mem_172_1_W0_addr),
    .W0_clk(mem_172_1_W0_clk),
    .W0_data(mem_172_1_W0_data),
    .W0_en(mem_172_1_W0_en),
    .W0_mask(mem_172_1_W0_mask)
  );
  split_mem_0_ext mem_172_2 (
    .R0_addr(mem_172_2_R0_addr),
    .R0_clk(mem_172_2_R0_clk),
    .R0_data(mem_172_2_R0_data),
    .R0_en(mem_172_2_R0_en),
    .W0_addr(mem_172_2_W0_addr),
    .W0_clk(mem_172_2_W0_clk),
    .W0_data(mem_172_2_W0_data),
    .W0_en(mem_172_2_W0_en),
    .W0_mask(mem_172_2_W0_mask)
  );
  split_mem_0_ext mem_172_3 (
    .R0_addr(mem_172_3_R0_addr),
    .R0_clk(mem_172_3_R0_clk),
    .R0_data(mem_172_3_R0_data),
    .R0_en(mem_172_3_R0_en),
    .W0_addr(mem_172_3_W0_addr),
    .W0_clk(mem_172_3_W0_clk),
    .W0_data(mem_172_3_W0_data),
    .W0_en(mem_172_3_W0_en),
    .W0_mask(mem_172_3_W0_mask)
  );
  split_mem_0_ext mem_172_4 (
    .R0_addr(mem_172_4_R0_addr),
    .R0_clk(mem_172_4_R0_clk),
    .R0_data(mem_172_4_R0_data),
    .R0_en(mem_172_4_R0_en),
    .W0_addr(mem_172_4_W0_addr),
    .W0_clk(mem_172_4_W0_clk),
    .W0_data(mem_172_4_W0_data),
    .W0_en(mem_172_4_W0_en),
    .W0_mask(mem_172_4_W0_mask)
  );
  split_mem_0_ext mem_172_5 (
    .R0_addr(mem_172_5_R0_addr),
    .R0_clk(mem_172_5_R0_clk),
    .R0_data(mem_172_5_R0_data),
    .R0_en(mem_172_5_R0_en),
    .W0_addr(mem_172_5_W0_addr),
    .W0_clk(mem_172_5_W0_clk),
    .W0_data(mem_172_5_W0_data),
    .W0_en(mem_172_5_W0_en),
    .W0_mask(mem_172_5_W0_mask)
  );
  split_mem_0_ext mem_172_6 (
    .R0_addr(mem_172_6_R0_addr),
    .R0_clk(mem_172_6_R0_clk),
    .R0_data(mem_172_6_R0_data),
    .R0_en(mem_172_6_R0_en),
    .W0_addr(mem_172_6_W0_addr),
    .W0_clk(mem_172_6_W0_clk),
    .W0_data(mem_172_6_W0_data),
    .W0_en(mem_172_6_W0_en),
    .W0_mask(mem_172_6_W0_mask)
  );
  split_mem_0_ext mem_172_7 (
    .R0_addr(mem_172_7_R0_addr),
    .R0_clk(mem_172_7_R0_clk),
    .R0_data(mem_172_7_R0_data),
    .R0_en(mem_172_7_R0_en),
    .W0_addr(mem_172_7_W0_addr),
    .W0_clk(mem_172_7_W0_clk),
    .W0_data(mem_172_7_W0_data),
    .W0_en(mem_172_7_W0_en),
    .W0_mask(mem_172_7_W0_mask)
  );
  split_mem_0_ext mem_173_0 (
    .R0_addr(mem_173_0_R0_addr),
    .R0_clk(mem_173_0_R0_clk),
    .R0_data(mem_173_0_R0_data),
    .R0_en(mem_173_0_R0_en),
    .W0_addr(mem_173_0_W0_addr),
    .W0_clk(mem_173_0_W0_clk),
    .W0_data(mem_173_0_W0_data),
    .W0_en(mem_173_0_W0_en),
    .W0_mask(mem_173_0_W0_mask)
  );
  split_mem_0_ext mem_173_1 (
    .R0_addr(mem_173_1_R0_addr),
    .R0_clk(mem_173_1_R0_clk),
    .R0_data(mem_173_1_R0_data),
    .R0_en(mem_173_1_R0_en),
    .W0_addr(mem_173_1_W0_addr),
    .W0_clk(mem_173_1_W0_clk),
    .W0_data(mem_173_1_W0_data),
    .W0_en(mem_173_1_W0_en),
    .W0_mask(mem_173_1_W0_mask)
  );
  split_mem_0_ext mem_173_2 (
    .R0_addr(mem_173_2_R0_addr),
    .R0_clk(mem_173_2_R0_clk),
    .R0_data(mem_173_2_R0_data),
    .R0_en(mem_173_2_R0_en),
    .W0_addr(mem_173_2_W0_addr),
    .W0_clk(mem_173_2_W0_clk),
    .W0_data(mem_173_2_W0_data),
    .W0_en(mem_173_2_W0_en),
    .W0_mask(mem_173_2_W0_mask)
  );
  split_mem_0_ext mem_173_3 (
    .R0_addr(mem_173_3_R0_addr),
    .R0_clk(mem_173_3_R0_clk),
    .R0_data(mem_173_3_R0_data),
    .R0_en(mem_173_3_R0_en),
    .W0_addr(mem_173_3_W0_addr),
    .W0_clk(mem_173_3_W0_clk),
    .W0_data(mem_173_3_W0_data),
    .W0_en(mem_173_3_W0_en),
    .W0_mask(mem_173_3_W0_mask)
  );
  split_mem_0_ext mem_173_4 (
    .R0_addr(mem_173_4_R0_addr),
    .R0_clk(mem_173_4_R0_clk),
    .R0_data(mem_173_4_R0_data),
    .R0_en(mem_173_4_R0_en),
    .W0_addr(mem_173_4_W0_addr),
    .W0_clk(mem_173_4_W0_clk),
    .W0_data(mem_173_4_W0_data),
    .W0_en(mem_173_4_W0_en),
    .W0_mask(mem_173_4_W0_mask)
  );
  split_mem_0_ext mem_173_5 (
    .R0_addr(mem_173_5_R0_addr),
    .R0_clk(mem_173_5_R0_clk),
    .R0_data(mem_173_5_R0_data),
    .R0_en(mem_173_5_R0_en),
    .W0_addr(mem_173_5_W0_addr),
    .W0_clk(mem_173_5_W0_clk),
    .W0_data(mem_173_5_W0_data),
    .W0_en(mem_173_5_W0_en),
    .W0_mask(mem_173_5_W0_mask)
  );
  split_mem_0_ext mem_173_6 (
    .R0_addr(mem_173_6_R0_addr),
    .R0_clk(mem_173_6_R0_clk),
    .R0_data(mem_173_6_R0_data),
    .R0_en(mem_173_6_R0_en),
    .W0_addr(mem_173_6_W0_addr),
    .W0_clk(mem_173_6_W0_clk),
    .W0_data(mem_173_6_W0_data),
    .W0_en(mem_173_6_W0_en),
    .W0_mask(mem_173_6_W0_mask)
  );
  split_mem_0_ext mem_173_7 (
    .R0_addr(mem_173_7_R0_addr),
    .R0_clk(mem_173_7_R0_clk),
    .R0_data(mem_173_7_R0_data),
    .R0_en(mem_173_7_R0_en),
    .W0_addr(mem_173_7_W0_addr),
    .W0_clk(mem_173_7_W0_clk),
    .W0_data(mem_173_7_W0_data),
    .W0_en(mem_173_7_W0_en),
    .W0_mask(mem_173_7_W0_mask)
  );
  split_mem_0_ext mem_174_0 (
    .R0_addr(mem_174_0_R0_addr),
    .R0_clk(mem_174_0_R0_clk),
    .R0_data(mem_174_0_R0_data),
    .R0_en(mem_174_0_R0_en),
    .W0_addr(mem_174_0_W0_addr),
    .W0_clk(mem_174_0_W0_clk),
    .W0_data(mem_174_0_W0_data),
    .W0_en(mem_174_0_W0_en),
    .W0_mask(mem_174_0_W0_mask)
  );
  split_mem_0_ext mem_174_1 (
    .R0_addr(mem_174_1_R0_addr),
    .R0_clk(mem_174_1_R0_clk),
    .R0_data(mem_174_1_R0_data),
    .R0_en(mem_174_1_R0_en),
    .W0_addr(mem_174_1_W0_addr),
    .W0_clk(mem_174_1_W0_clk),
    .W0_data(mem_174_1_W0_data),
    .W0_en(mem_174_1_W0_en),
    .W0_mask(mem_174_1_W0_mask)
  );
  split_mem_0_ext mem_174_2 (
    .R0_addr(mem_174_2_R0_addr),
    .R0_clk(mem_174_2_R0_clk),
    .R0_data(mem_174_2_R0_data),
    .R0_en(mem_174_2_R0_en),
    .W0_addr(mem_174_2_W0_addr),
    .W0_clk(mem_174_2_W0_clk),
    .W0_data(mem_174_2_W0_data),
    .W0_en(mem_174_2_W0_en),
    .W0_mask(mem_174_2_W0_mask)
  );
  split_mem_0_ext mem_174_3 (
    .R0_addr(mem_174_3_R0_addr),
    .R0_clk(mem_174_3_R0_clk),
    .R0_data(mem_174_3_R0_data),
    .R0_en(mem_174_3_R0_en),
    .W0_addr(mem_174_3_W0_addr),
    .W0_clk(mem_174_3_W0_clk),
    .W0_data(mem_174_3_W0_data),
    .W0_en(mem_174_3_W0_en),
    .W0_mask(mem_174_3_W0_mask)
  );
  split_mem_0_ext mem_174_4 (
    .R0_addr(mem_174_4_R0_addr),
    .R0_clk(mem_174_4_R0_clk),
    .R0_data(mem_174_4_R0_data),
    .R0_en(mem_174_4_R0_en),
    .W0_addr(mem_174_4_W0_addr),
    .W0_clk(mem_174_4_W0_clk),
    .W0_data(mem_174_4_W0_data),
    .W0_en(mem_174_4_W0_en),
    .W0_mask(mem_174_4_W0_mask)
  );
  split_mem_0_ext mem_174_5 (
    .R0_addr(mem_174_5_R0_addr),
    .R0_clk(mem_174_5_R0_clk),
    .R0_data(mem_174_5_R0_data),
    .R0_en(mem_174_5_R0_en),
    .W0_addr(mem_174_5_W0_addr),
    .W0_clk(mem_174_5_W0_clk),
    .W0_data(mem_174_5_W0_data),
    .W0_en(mem_174_5_W0_en),
    .W0_mask(mem_174_5_W0_mask)
  );
  split_mem_0_ext mem_174_6 (
    .R0_addr(mem_174_6_R0_addr),
    .R0_clk(mem_174_6_R0_clk),
    .R0_data(mem_174_6_R0_data),
    .R0_en(mem_174_6_R0_en),
    .W0_addr(mem_174_6_W0_addr),
    .W0_clk(mem_174_6_W0_clk),
    .W0_data(mem_174_6_W0_data),
    .W0_en(mem_174_6_W0_en),
    .W0_mask(mem_174_6_W0_mask)
  );
  split_mem_0_ext mem_174_7 (
    .R0_addr(mem_174_7_R0_addr),
    .R0_clk(mem_174_7_R0_clk),
    .R0_data(mem_174_7_R0_data),
    .R0_en(mem_174_7_R0_en),
    .W0_addr(mem_174_7_W0_addr),
    .W0_clk(mem_174_7_W0_clk),
    .W0_data(mem_174_7_W0_data),
    .W0_en(mem_174_7_W0_en),
    .W0_mask(mem_174_7_W0_mask)
  );
  split_mem_0_ext mem_175_0 (
    .R0_addr(mem_175_0_R0_addr),
    .R0_clk(mem_175_0_R0_clk),
    .R0_data(mem_175_0_R0_data),
    .R0_en(mem_175_0_R0_en),
    .W0_addr(mem_175_0_W0_addr),
    .W0_clk(mem_175_0_W0_clk),
    .W0_data(mem_175_0_W0_data),
    .W0_en(mem_175_0_W0_en),
    .W0_mask(mem_175_0_W0_mask)
  );
  split_mem_0_ext mem_175_1 (
    .R0_addr(mem_175_1_R0_addr),
    .R0_clk(mem_175_1_R0_clk),
    .R0_data(mem_175_1_R0_data),
    .R0_en(mem_175_1_R0_en),
    .W0_addr(mem_175_1_W0_addr),
    .W0_clk(mem_175_1_W0_clk),
    .W0_data(mem_175_1_W0_data),
    .W0_en(mem_175_1_W0_en),
    .W0_mask(mem_175_1_W0_mask)
  );
  split_mem_0_ext mem_175_2 (
    .R0_addr(mem_175_2_R0_addr),
    .R0_clk(mem_175_2_R0_clk),
    .R0_data(mem_175_2_R0_data),
    .R0_en(mem_175_2_R0_en),
    .W0_addr(mem_175_2_W0_addr),
    .W0_clk(mem_175_2_W0_clk),
    .W0_data(mem_175_2_W0_data),
    .W0_en(mem_175_2_W0_en),
    .W0_mask(mem_175_2_W0_mask)
  );
  split_mem_0_ext mem_175_3 (
    .R0_addr(mem_175_3_R0_addr),
    .R0_clk(mem_175_3_R0_clk),
    .R0_data(mem_175_3_R0_data),
    .R0_en(mem_175_3_R0_en),
    .W0_addr(mem_175_3_W0_addr),
    .W0_clk(mem_175_3_W0_clk),
    .W0_data(mem_175_3_W0_data),
    .W0_en(mem_175_3_W0_en),
    .W0_mask(mem_175_3_W0_mask)
  );
  split_mem_0_ext mem_175_4 (
    .R0_addr(mem_175_4_R0_addr),
    .R0_clk(mem_175_4_R0_clk),
    .R0_data(mem_175_4_R0_data),
    .R0_en(mem_175_4_R0_en),
    .W0_addr(mem_175_4_W0_addr),
    .W0_clk(mem_175_4_W0_clk),
    .W0_data(mem_175_4_W0_data),
    .W0_en(mem_175_4_W0_en),
    .W0_mask(mem_175_4_W0_mask)
  );
  split_mem_0_ext mem_175_5 (
    .R0_addr(mem_175_5_R0_addr),
    .R0_clk(mem_175_5_R0_clk),
    .R0_data(mem_175_5_R0_data),
    .R0_en(mem_175_5_R0_en),
    .W0_addr(mem_175_5_W0_addr),
    .W0_clk(mem_175_5_W0_clk),
    .W0_data(mem_175_5_W0_data),
    .W0_en(mem_175_5_W0_en),
    .W0_mask(mem_175_5_W0_mask)
  );
  split_mem_0_ext mem_175_6 (
    .R0_addr(mem_175_6_R0_addr),
    .R0_clk(mem_175_6_R0_clk),
    .R0_data(mem_175_6_R0_data),
    .R0_en(mem_175_6_R0_en),
    .W0_addr(mem_175_6_W0_addr),
    .W0_clk(mem_175_6_W0_clk),
    .W0_data(mem_175_6_W0_data),
    .W0_en(mem_175_6_W0_en),
    .W0_mask(mem_175_6_W0_mask)
  );
  split_mem_0_ext mem_175_7 (
    .R0_addr(mem_175_7_R0_addr),
    .R0_clk(mem_175_7_R0_clk),
    .R0_data(mem_175_7_R0_data),
    .R0_en(mem_175_7_R0_en),
    .W0_addr(mem_175_7_W0_addr),
    .W0_clk(mem_175_7_W0_clk),
    .W0_data(mem_175_7_W0_data),
    .W0_en(mem_175_7_W0_en),
    .W0_mask(mem_175_7_W0_mask)
  );
  split_mem_0_ext mem_176_0 (
    .R0_addr(mem_176_0_R0_addr),
    .R0_clk(mem_176_0_R0_clk),
    .R0_data(mem_176_0_R0_data),
    .R0_en(mem_176_0_R0_en),
    .W0_addr(mem_176_0_W0_addr),
    .W0_clk(mem_176_0_W0_clk),
    .W0_data(mem_176_0_W0_data),
    .W0_en(mem_176_0_W0_en),
    .W0_mask(mem_176_0_W0_mask)
  );
  split_mem_0_ext mem_176_1 (
    .R0_addr(mem_176_1_R0_addr),
    .R0_clk(mem_176_1_R0_clk),
    .R0_data(mem_176_1_R0_data),
    .R0_en(mem_176_1_R0_en),
    .W0_addr(mem_176_1_W0_addr),
    .W0_clk(mem_176_1_W0_clk),
    .W0_data(mem_176_1_W0_data),
    .W0_en(mem_176_1_W0_en),
    .W0_mask(mem_176_1_W0_mask)
  );
  split_mem_0_ext mem_176_2 (
    .R0_addr(mem_176_2_R0_addr),
    .R0_clk(mem_176_2_R0_clk),
    .R0_data(mem_176_2_R0_data),
    .R0_en(mem_176_2_R0_en),
    .W0_addr(mem_176_2_W0_addr),
    .W0_clk(mem_176_2_W0_clk),
    .W0_data(mem_176_2_W0_data),
    .W0_en(mem_176_2_W0_en),
    .W0_mask(mem_176_2_W0_mask)
  );
  split_mem_0_ext mem_176_3 (
    .R0_addr(mem_176_3_R0_addr),
    .R0_clk(mem_176_3_R0_clk),
    .R0_data(mem_176_3_R0_data),
    .R0_en(mem_176_3_R0_en),
    .W0_addr(mem_176_3_W0_addr),
    .W0_clk(mem_176_3_W0_clk),
    .W0_data(mem_176_3_W0_data),
    .W0_en(mem_176_3_W0_en),
    .W0_mask(mem_176_3_W0_mask)
  );
  split_mem_0_ext mem_176_4 (
    .R0_addr(mem_176_4_R0_addr),
    .R0_clk(mem_176_4_R0_clk),
    .R0_data(mem_176_4_R0_data),
    .R0_en(mem_176_4_R0_en),
    .W0_addr(mem_176_4_W0_addr),
    .W0_clk(mem_176_4_W0_clk),
    .W0_data(mem_176_4_W0_data),
    .W0_en(mem_176_4_W0_en),
    .W0_mask(mem_176_4_W0_mask)
  );
  split_mem_0_ext mem_176_5 (
    .R0_addr(mem_176_5_R0_addr),
    .R0_clk(mem_176_5_R0_clk),
    .R0_data(mem_176_5_R0_data),
    .R0_en(mem_176_5_R0_en),
    .W0_addr(mem_176_5_W0_addr),
    .W0_clk(mem_176_5_W0_clk),
    .W0_data(mem_176_5_W0_data),
    .W0_en(mem_176_5_W0_en),
    .W0_mask(mem_176_5_W0_mask)
  );
  split_mem_0_ext mem_176_6 (
    .R0_addr(mem_176_6_R0_addr),
    .R0_clk(mem_176_6_R0_clk),
    .R0_data(mem_176_6_R0_data),
    .R0_en(mem_176_6_R0_en),
    .W0_addr(mem_176_6_W0_addr),
    .W0_clk(mem_176_6_W0_clk),
    .W0_data(mem_176_6_W0_data),
    .W0_en(mem_176_6_W0_en),
    .W0_mask(mem_176_6_W0_mask)
  );
  split_mem_0_ext mem_176_7 (
    .R0_addr(mem_176_7_R0_addr),
    .R0_clk(mem_176_7_R0_clk),
    .R0_data(mem_176_7_R0_data),
    .R0_en(mem_176_7_R0_en),
    .W0_addr(mem_176_7_W0_addr),
    .W0_clk(mem_176_7_W0_clk),
    .W0_data(mem_176_7_W0_data),
    .W0_en(mem_176_7_W0_en),
    .W0_mask(mem_176_7_W0_mask)
  );
  split_mem_0_ext mem_177_0 (
    .R0_addr(mem_177_0_R0_addr),
    .R0_clk(mem_177_0_R0_clk),
    .R0_data(mem_177_0_R0_data),
    .R0_en(mem_177_0_R0_en),
    .W0_addr(mem_177_0_W0_addr),
    .W0_clk(mem_177_0_W0_clk),
    .W0_data(mem_177_0_W0_data),
    .W0_en(mem_177_0_W0_en),
    .W0_mask(mem_177_0_W0_mask)
  );
  split_mem_0_ext mem_177_1 (
    .R0_addr(mem_177_1_R0_addr),
    .R0_clk(mem_177_1_R0_clk),
    .R0_data(mem_177_1_R0_data),
    .R0_en(mem_177_1_R0_en),
    .W0_addr(mem_177_1_W0_addr),
    .W0_clk(mem_177_1_W0_clk),
    .W0_data(mem_177_1_W0_data),
    .W0_en(mem_177_1_W0_en),
    .W0_mask(mem_177_1_W0_mask)
  );
  split_mem_0_ext mem_177_2 (
    .R0_addr(mem_177_2_R0_addr),
    .R0_clk(mem_177_2_R0_clk),
    .R0_data(mem_177_2_R0_data),
    .R0_en(mem_177_2_R0_en),
    .W0_addr(mem_177_2_W0_addr),
    .W0_clk(mem_177_2_W0_clk),
    .W0_data(mem_177_2_W0_data),
    .W0_en(mem_177_2_W0_en),
    .W0_mask(mem_177_2_W0_mask)
  );
  split_mem_0_ext mem_177_3 (
    .R0_addr(mem_177_3_R0_addr),
    .R0_clk(mem_177_3_R0_clk),
    .R0_data(mem_177_3_R0_data),
    .R0_en(mem_177_3_R0_en),
    .W0_addr(mem_177_3_W0_addr),
    .W0_clk(mem_177_3_W0_clk),
    .W0_data(mem_177_3_W0_data),
    .W0_en(mem_177_3_W0_en),
    .W0_mask(mem_177_3_W0_mask)
  );
  split_mem_0_ext mem_177_4 (
    .R0_addr(mem_177_4_R0_addr),
    .R0_clk(mem_177_4_R0_clk),
    .R0_data(mem_177_4_R0_data),
    .R0_en(mem_177_4_R0_en),
    .W0_addr(mem_177_4_W0_addr),
    .W0_clk(mem_177_4_W0_clk),
    .W0_data(mem_177_4_W0_data),
    .W0_en(mem_177_4_W0_en),
    .W0_mask(mem_177_4_W0_mask)
  );
  split_mem_0_ext mem_177_5 (
    .R0_addr(mem_177_5_R0_addr),
    .R0_clk(mem_177_5_R0_clk),
    .R0_data(mem_177_5_R0_data),
    .R0_en(mem_177_5_R0_en),
    .W0_addr(mem_177_5_W0_addr),
    .W0_clk(mem_177_5_W0_clk),
    .W0_data(mem_177_5_W0_data),
    .W0_en(mem_177_5_W0_en),
    .W0_mask(mem_177_5_W0_mask)
  );
  split_mem_0_ext mem_177_6 (
    .R0_addr(mem_177_6_R0_addr),
    .R0_clk(mem_177_6_R0_clk),
    .R0_data(mem_177_6_R0_data),
    .R0_en(mem_177_6_R0_en),
    .W0_addr(mem_177_6_W0_addr),
    .W0_clk(mem_177_6_W0_clk),
    .W0_data(mem_177_6_W0_data),
    .W0_en(mem_177_6_W0_en),
    .W0_mask(mem_177_6_W0_mask)
  );
  split_mem_0_ext mem_177_7 (
    .R0_addr(mem_177_7_R0_addr),
    .R0_clk(mem_177_7_R0_clk),
    .R0_data(mem_177_7_R0_data),
    .R0_en(mem_177_7_R0_en),
    .W0_addr(mem_177_7_W0_addr),
    .W0_clk(mem_177_7_W0_clk),
    .W0_data(mem_177_7_W0_data),
    .W0_en(mem_177_7_W0_en),
    .W0_mask(mem_177_7_W0_mask)
  );
  split_mem_0_ext mem_178_0 (
    .R0_addr(mem_178_0_R0_addr),
    .R0_clk(mem_178_0_R0_clk),
    .R0_data(mem_178_0_R0_data),
    .R0_en(mem_178_0_R0_en),
    .W0_addr(mem_178_0_W0_addr),
    .W0_clk(mem_178_0_W0_clk),
    .W0_data(mem_178_0_W0_data),
    .W0_en(mem_178_0_W0_en),
    .W0_mask(mem_178_0_W0_mask)
  );
  split_mem_0_ext mem_178_1 (
    .R0_addr(mem_178_1_R0_addr),
    .R0_clk(mem_178_1_R0_clk),
    .R0_data(mem_178_1_R0_data),
    .R0_en(mem_178_1_R0_en),
    .W0_addr(mem_178_1_W0_addr),
    .W0_clk(mem_178_1_W0_clk),
    .W0_data(mem_178_1_W0_data),
    .W0_en(mem_178_1_W0_en),
    .W0_mask(mem_178_1_W0_mask)
  );
  split_mem_0_ext mem_178_2 (
    .R0_addr(mem_178_2_R0_addr),
    .R0_clk(mem_178_2_R0_clk),
    .R0_data(mem_178_2_R0_data),
    .R0_en(mem_178_2_R0_en),
    .W0_addr(mem_178_2_W0_addr),
    .W0_clk(mem_178_2_W0_clk),
    .W0_data(mem_178_2_W0_data),
    .W0_en(mem_178_2_W0_en),
    .W0_mask(mem_178_2_W0_mask)
  );
  split_mem_0_ext mem_178_3 (
    .R0_addr(mem_178_3_R0_addr),
    .R0_clk(mem_178_3_R0_clk),
    .R0_data(mem_178_3_R0_data),
    .R0_en(mem_178_3_R0_en),
    .W0_addr(mem_178_3_W0_addr),
    .W0_clk(mem_178_3_W0_clk),
    .W0_data(mem_178_3_W0_data),
    .W0_en(mem_178_3_W0_en),
    .W0_mask(mem_178_3_W0_mask)
  );
  split_mem_0_ext mem_178_4 (
    .R0_addr(mem_178_4_R0_addr),
    .R0_clk(mem_178_4_R0_clk),
    .R0_data(mem_178_4_R0_data),
    .R0_en(mem_178_4_R0_en),
    .W0_addr(mem_178_4_W0_addr),
    .W0_clk(mem_178_4_W0_clk),
    .W0_data(mem_178_4_W0_data),
    .W0_en(mem_178_4_W0_en),
    .W0_mask(mem_178_4_W0_mask)
  );
  split_mem_0_ext mem_178_5 (
    .R0_addr(mem_178_5_R0_addr),
    .R0_clk(mem_178_5_R0_clk),
    .R0_data(mem_178_5_R0_data),
    .R0_en(mem_178_5_R0_en),
    .W0_addr(mem_178_5_W0_addr),
    .W0_clk(mem_178_5_W0_clk),
    .W0_data(mem_178_5_W0_data),
    .W0_en(mem_178_5_W0_en),
    .W0_mask(mem_178_5_W0_mask)
  );
  split_mem_0_ext mem_178_6 (
    .R0_addr(mem_178_6_R0_addr),
    .R0_clk(mem_178_6_R0_clk),
    .R0_data(mem_178_6_R0_data),
    .R0_en(mem_178_6_R0_en),
    .W0_addr(mem_178_6_W0_addr),
    .W0_clk(mem_178_6_W0_clk),
    .W0_data(mem_178_6_W0_data),
    .W0_en(mem_178_6_W0_en),
    .W0_mask(mem_178_6_W0_mask)
  );
  split_mem_0_ext mem_178_7 (
    .R0_addr(mem_178_7_R0_addr),
    .R0_clk(mem_178_7_R0_clk),
    .R0_data(mem_178_7_R0_data),
    .R0_en(mem_178_7_R0_en),
    .W0_addr(mem_178_7_W0_addr),
    .W0_clk(mem_178_7_W0_clk),
    .W0_data(mem_178_7_W0_data),
    .W0_en(mem_178_7_W0_en),
    .W0_mask(mem_178_7_W0_mask)
  );
  split_mem_0_ext mem_179_0 (
    .R0_addr(mem_179_0_R0_addr),
    .R0_clk(mem_179_0_R0_clk),
    .R0_data(mem_179_0_R0_data),
    .R0_en(mem_179_0_R0_en),
    .W0_addr(mem_179_0_W0_addr),
    .W0_clk(mem_179_0_W0_clk),
    .W0_data(mem_179_0_W0_data),
    .W0_en(mem_179_0_W0_en),
    .W0_mask(mem_179_0_W0_mask)
  );
  split_mem_0_ext mem_179_1 (
    .R0_addr(mem_179_1_R0_addr),
    .R0_clk(mem_179_1_R0_clk),
    .R0_data(mem_179_1_R0_data),
    .R0_en(mem_179_1_R0_en),
    .W0_addr(mem_179_1_W0_addr),
    .W0_clk(mem_179_1_W0_clk),
    .W0_data(mem_179_1_W0_data),
    .W0_en(mem_179_1_W0_en),
    .W0_mask(mem_179_1_W0_mask)
  );
  split_mem_0_ext mem_179_2 (
    .R0_addr(mem_179_2_R0_addr),
    .R0_clk(mem_179_2_R0_clk),
    .R0_data(mem_179_2_R0_data),
    .R0_en(mem_179_2_R0_en),
    .W0_addr(mem_179_2_W0_addr),
    .W0_clk(mem_179_2_W0_clk),
    .W0_data(mem_179_2_W0_data),
    .W0_en(mem_179_2_W0_en),
    .W0_mask(mem_179_2_W0_mask)
  );
  split_mem_0_ext mem_179_3 (
    .R0_addr(mem_179_3_R0_addr),
    .R0_clk(mem_179_3_R0_clk),
    .R0_data(mem_179_3_R0_data),
    .R0_en(mem_179_3_R0_en),
    .W0_addr(mem_179_3_W0_addr),
    .W0_clk(mem_179_3_W0_clk),
    .W0_data(mem_179_3_W0_data),
    .W0_en(mem_179_3_W0_en),
    .W0_mask(mem_179_3_W0_mask)
  );
  split_mem_0_ext mem_179_4 (
    .R0_addr(mem_179_4_R0_addr),
    .R0_clk(mem_179_4_R0_clk),
    .R0_data(mem_179_4_R0_data),
    .R0_en(mem_179_4_R0_en),
    .W0_addr(mem_179_4_W0_addr),
    .W0_clk(mem_179_4_W0_clk),
    .W0_data(mem_179_4_W0_data),
    .W0_en(mem_179_4_W0_en),
    .W0_mask(mem_179_4_W0_mask)
  );
  split_mem_0_ext mem_179_5 (
    .R0_addr(mem_179_5_R0_addr),
    .R0_clk(mem_179_5_R0_clk),
    .R0_data(mem_179_5_R0_data),
    .R0_en(mem_179_5_R0_en),
    .W0_addr(mem_179_5_W0_addr),
    .W0_clk(mem_179_5_W0_clk),
    .W0_data(mem_179_5_W0_data),
    .W0_en(mem_179_5_W0_en),
    .W0_mask(mem_179_5_W0_mask)
  );
  split_mem_0_ext mem_179_6 (
    .R0_addr(mem_179_6_R0_addr),
    .R0_clk(mem_179_6_R0_clk),
    .R0_data(mem_179_6_R0_data),
    .R0_en(mem_179_6_R0_en),
    .W0_addr(mem_179_6_W0_addr),
    .W0_clk(mem_179_6_W0_clk),
    .W0_data(mem_179_6_W0_data),
    .W0_en(mem_179_6_W0_en),
    .W0_mask(mem_179_6_W0_mask)
  );
  split_mem_0_ext mem_179_7 (
    .R0_addr(mem_179_7_R0_addr),
    .R0_clk(mem_179_7_R0_clk),
    .R0_data(mem_179_7_R0_data),
    .R0_en(mem_179_7_R0_en),
    .W0_addr(mem_179_7_W0_addr),
    .W0_clk(mem_179_7_W0_clk),
    .W0_data(mem_179_7_W0_data),
    .W0_en(mem_179_7_W0_en),
    .W0_mask(mem_179_7_W0_mask)
  );
  split_mem_0_ext mem_180_0 (
    .R0_addr(mem_180_0_R0_addr),
    .R0_clk(mem_180_0_R0_clk),
    .R0_data(mem_180_0_R0_data),
    .R0_en(mem_180_0_R0_en),
    .W0_addr(mem_180_0_W0_addr),
    .W0_clk(mem_180_0_W0_clk),
    .W0_data(mem_180_0_W0_data),
    .W0_en(mem_180_0_W0_en),
    .W0_mask(mem_180_0_W0_mask)
  );
  split_mem_0_ext mem_180_1 (
    .R0_addr(mem_180_1_R0_addr),
    .R0_clk(mem_180_1_R0_clk),
    .R0_data(mem_180_1_R0_data),
    .R0_en(mem_180_1_R0_en),
    .W0_addr(mem_180_1_W0_addr),
    .W0_clk(mem_180_1_W0_clk),
    .W0_data(mem_180_1_W0_data),
    .W0_en(mem_180_1_W0_en),
    .W0_mask(mem_180_1_W0_mask)
  );
  split_mem_0_ext mem_180_2 (
    .R0_addr(mem_180_2_R0_addr),
    .R0_clk(mem_180_2_R0_clk),
    .R0_data(mem_180_2_R0_data),
    .R0_en(mem_180_2_R0_en),
    .W0_addr(mem_180_2_W0_addr),
    .W0_clk(mem_180_2_W0_clk),
    .W0_data(mem_180_2_W0_data),
    .W0_en(mem_180_2_W0_en),
    .W0_mask(mem_180_2_W0_mask)
  );
  split_mem_0_ext mem_180_3 (
    .R0_addr(mem_180_3_R0_addr),
    .R0_clk(mem_180_3_R0_clk),
    .R0_data(mem_180_3_R0_data),
    .R0_en(mem_180_3_R0_en),
    .W0_addr(mem_180_3_W0_addr),
    .W0_clk(mem_180_3_W0_clk),
    .W0_data(mem_180_3_W0_data),
    .W0_en(mem_180_3_W0_en),
    .W0_mask(mem_180_3_W0_mask)
  );
  split_mem_0_ext mem_180_4 (
    .R0_addr(mem_180_4_R0_addr),
    .R0_clk(mem_180_4_R0_clk),
    .R0_data(mem_180_4_R0_data),
    .R0_en(mem_180_4_R0_en),
    .W0_addr(mem_180_4_W0_addr),
    .W0_clk(mem_180_4_W0_clk),
    .W0_data(mem_180_4_W0_data),
    .W0_en(mem_180_4_W0_en),
    .W0_mask(mem_180_4_W0_mask)
  );
  split_mem_0_ext mem_180_5 (
    .R0_addr(mem_180_5_R0_addr),
    .R0_clk(mem_180_5_R0_clk),
    .R0_data(mem_180_5_R0_data),
    .R0_en(mem_180_5_R0_en),
    .W0_addr(mem_180_5_W0_addr),
    .W0_clk(mem_180_5_W0_clk),
    .W0_data(mem_180_5_W0_data),
    .W0_en(mem_180_5_W0_en),
    .W0_mask(mem_180_5_W0_mask)
  );
  split_mem_0_ext mem_180_6 (
    .R0_addr(mem_180_6_R0_addr),
    .R0_clk(mem_180_6_R0_clk),
    .R0_data(mem_180_6_R0_data),
    .R0_en(mem_180_6_R0_en),
    .W0_addr(mem_180_6_W0_addr),
    .W0_clk(mem_180_6_W0_clk),
    .W0_data(mem_180_6_W0_data),
    .W0_en(mem_180_6_W0_en),
    .W0_mask(mem_180_6_W0_mask)
  );
  split_mem_0_ext mem_180_7 (
    .R0_addr(mem_180_7_R0_addr),
    .R0_clk(mem_180_7_R0_clk),
    .R0_data(mem_180_7_R0_data),
    .R0_en(mem_180_7_R0_en),
    .W0_addr(mem_180_7_W0_addr),
    .W0_clk(mem_180_7_W0_clk),
    .W0_data(mem_180_7_W0_data),
    .W0_en(mem_180_7_W0_en),
    .W0_mask(mem_180_7_W0_mask)
  );
  split_mem_0_ext mem_181_0 (
    .R0_addr(mem_181_0_R0_addr),
    .R0_clk(mem_181_0_R0_clk),
    .R0_data(mem_181_0_R0_data),
    .R0_en(mem_181_0_R0_en),
    .W0_addr(mem_181_0_W0_addr),
    .W0_clk(mem_181_0_W0_clk),
    .W0_data(mem_181_0_W0_data),
    .W0_en(mem_181_0_W0_en),
    .W0_mask(mem_181_0_W0_mask)
  );
  split_mem_0_ext mem_181_1 (
    .R0_addr(mem_181_1_R0_addr),
    .R0_clk(mem_181_1_R0_clk),
    .R0_data(mem_181_1_R0_data),
    .R0_en(mem_181_1_R0_en),
    .W0_addr(mem_181_1_W0_addr),
    .W0_clk(mem_181_1_W0_clk),
    .W0_data(mem_181_1_W0_data),
    .W0_en(mem_181_1_W0_en),
    .W0_mask(mem_181_1_W0_mask)
  );
  split_mem_0_ext mem_181_2 (
    .R0_addr(mem_181_2_R0_addr),
    .R0_clk(mem_181_2_R0_clk),
    .R0_data(mem_181_2_R0_data),
    .R0_en(mem_181_2_R0_en),
    .W0_addr(mem_181_2_W0_addr),
    .W0_clk(mem_181_2_W0_clk),
    .W0_data(mem_181_2_W0_data),
    .W0_en(mem_181_2_W0_en),
    .W0_mask(mem_181_2_W0_mask)
  );
  split_mem_0_ext mem_181_3 (
    .R0_addr(mem_181_3_R0_addr),
    .R0_clk(mem_181_3_R0_clk),
    .R0_data(mem_181_3_R0_data),
    .R0_en(mem_181_3_R0_en),
    .W0_addr(mem_181_3_W0_addr),
    .W0_clk(mem_181_3_W0_clk),
    .W0_data(mem_181_3_W0_data),
    .W0_en(mem_181_3_W0_en),
    .W0_mask(mem_181_3_W0_mask)
  );
  split_mem_0_ext mem_181_4 (
    .R0_addr(mem_181_4_R0_addr),
    .R0_clk(mem_181_4_R0_clk),
    .R0_data(mem_181_4_R0_data),
    .R0_en(mem_181_4_R0_en),
    .W0_addr(mem_181_4_W0_addr),
    .W0_clk(mem_181_4_W0_clk),
    .W0_data(mem_181_4_W0_data),
    .W0_en(mem_181_4_W0_en),
    .W0_mask(mem_181_4_W0_mask)
  );
  split_mem_0_ext mem_181_5 (
    .R0_addr(mem_181_5_R0_addr),
    .R0_clk(mem_181_5_R0_clk),
    .R0_data(mem_181_5_R0_data),
    .R0_en(mem_181_5_R0_en),
    .W0_addr(mem_181_5_W0_addr),
    .W0_clk(mem_181_5_W0_clk),
    .W0_data(mem_181_5_W0_data),
    .W0_en(mem_181_5_W0_en),
    .W0_mask(mem_181_5_W0_mask)
  );
  split_mem_0_ext mem_181_6 (
    .R0_addr(mem_181_6_R0_addr),
    .R0_clk(mem_181_6_R0_clk),
    .R0_data(mem_181_6_R0_data),
    .R0_en(mem_181_6_R0_en),
    .W0_addr(mem_181_6_W0_addr),
    .W0_clk(mem_181_6_W0_clk),
    .W0_data(mem_181_6_W0_data),
    .W0_en(mem_181_6_W0_en),
    .W0_mask(mem_181_6_W0_mask)
  );
  split_mem_0_ext mem_181_7 (
    .R0_addr(mem_181_7_R0_addr),
    .R0_clk(mem_181_7_R0_clk),
    .R0_data(mem_181_7_R0_data),
    .R0_en(mem_181_7_R0_en),
    .W0_addr(mem_181_7_W0_addr),
    .W0_clk(mem_181_7_W0_clk),
    .W0_data(mem_181_7_W0_data),
    .W0_en(mem_181_7_W0_en),
    .W0_mask(mem_181_7_W0_mask)
  );
  split_mem_0_ext mem_182_0 (
    .R0_addr(mem_182_0_R0_addr),
    .R0_clk(mem_182_0_R0_clk),
    .R0_data(mem_182_0_R0_data),
    .R0_en(mem_182_0_R0_en),
    .W0_addr(mem_182_0_W0_addr),
    .W0_clk(mem_182_0_W0_clk),
    .W0_data(mem_182_0_W0_data),
    .W0_en(mem_182_0_W0_en),
    .W0_mask(mem_182_0_W0_mask)
  );
  split_mem_0_ext mem_182_1 (
    .R0_addr(mem_182_1_R0_addr),
    .R0_clk(mem_182_1_R0_clk),
    .R0_data(mem_182_1_R0_data),
    .R0_en(mem_182_1_R0_en),
    .W0_addr(mem_182_1_W0_addr),
    .W0_clk(mem_182_1_W0_clk),
    .W0_data(mem_182_1_W0_data),
    .W0_en(mem_182_1_W0_en),
    .W0_mask(mem_182_1_W0_mask)
  );
  split_mem_0_ext mem_182_2 (
    .R0_addr(mem_182_2_R0_addr),
    .R0_clk(mem_182_2_R0_clk),
    .R0_data(mem_182_2_R0_data),
    .R0_en(mem_182_2_R0_en),
    .W0_addr(mem_182_2_W0_addr),
    .W0_clk(mem_182_2_W0_clk),
    .W0_data(mem_182_2_W0_data),
    .W0_en(mem_182_2_W0_en),
    .W0_mask(mem_182_2_W0_mask)
  );
  split_mem_0_ext mem_182_3 (
    .R0_addr(mem_182_3_R0_addr),
    .R0_clk(mem_182_3_R0_clk),
    .R0_data(mem_182_3_R0_data),
    .R0_en(mem_182_3_R0_en),
    .W0_addr(mem_182_3_W0_addr),
    .W0_clk(mem_182_3_W0_clk),
    .W0_data(mem_182_3_W0_data),
    .W0_en(mem_182_3_W0_en),
    .W0_mask(mem_182_3_W0_mask)
  );
  split_mem_0_ext mem_182_4 (
    .R0_addr(mem_182_4_R0_addr),
    .R0_clk(mem_182_4_R0_clk),
    .R0_data(mem_182_4_R0_data),
    .R0_en(mem_182_4_R0_en),
    .W0_addr(mem_182_4_W0_addr),
    .W0_clk(mem_182_4_W0_clk),
    .W0_data(mem_182_4_W0_data),
    .W0_en(mem_182_4_W0_en),
    .W0_mask(mem_182_4_W0_mask)
  );
  split_mem_0_ext mem_182_5 (
    .R0_addr(mem_182_5_R0_addr),
    .R0_clk(mem_182_5_R0_clk),
    .R0_data(mem_182_5_R0_data),
    .R0_en(mem_182_5_R0_en),
    .W0_addr(mem_182_5_W0_addr),
    .W0_clk(mem_182_5_W0_clk),
    .W0_data(mem_182_5_W0_data),
    .W0_en(mem_182_5_W0_en),
    .W0_mask(mem_182_5_W0_mask)
  );
  split_mem_0_ext mem_182_6 (
    .R0_addr(mem_182_6_R0_addr),
    .R0_clk(mem_182_6_R0_clk),
    .R0_data(mem_182_6_R0_data),
    .R0_en(mem_182_6_R0_en),
    .W0_addr(mem_182_6_W0_addr),
    .W0_clk(mem_182_6_W0_clk),
    .W0_data(mem_182_6_W0_data),
    .W0_en(mem_182_6_W0_en),
    .W0_mask(mem_182_6_W0_mask)
  );
  split_mem_0_ext mem_182_7 (
    .R0_addr(mem_182_7_R0_addr),
    .R0_clk(mem_182_7_R0_clk),
    .R0_data(mem_182_7_R0_data),
    .R0_en(mem_182_7_R0_en),
    .W0_addr(mem_182_7_W0_addr),
    .W0_clk(mem_182_7_W0_clk),
    .W0_data(mem_182_7_W0_data),
    .W0_en(mem_182_7_W0_en),
    .W0_mask(mem_182_7_W0_mask)
  );
  split_mem_0_ext mem_183_0 (
    .R0_addr(mem_183_0_R0_addr),
    .R0_clk(mem_183_0_R0_clk),
    .R0_data(mem_183_0_R0_data),
    .R0_en(mem_183_0_R0_en),
    .W0_addr(mem_183_0_W0_addr),
    .W0_clk(mem_183_0_W0_clk),
    .W0_data(mem_183_0_W0_data),
    .W0_en(mem_183_0_W0_en),
    .W0_mask(mem_183_0_W0_mask)
  );
  split_mem_0_ext mem_183_1 (
    .R0_addr(mem_183_1_R0_addr),
    .R0_clk(mem_183_1_R0_clk),
    .R0_data(mem_183_1_R0_data),
    .R0_en(mem_183_1_R0_en),
    .W0_addr(mem_183_1_W0_addr),
    .W0_clk(mem_183_1_W0_clk),
    .W0_data(mem_183_1_W0_data),
    .W0_en(mem_183_1_W0_en),
    .W0_mask(mem_183_1_W0_mask)
  );
  split_mem_0_ext mem_183_2 (
    .R0_addr(mem_183_2_R0_addr),
    .R0_clk(mem_183_2_R0_clk),
    .R0_data(mem_183_2_R0_data),
    .R0_en(mem_183_2_R0_en),
    .W0_addr(mem_183_2_W0_addr),
    .W0_clk(mem_183_2_W0_clk),
    .W0_data(mem_183_2_W0_data),
    .W0_en(mem_183_2_W0_en),
    .W0_mask(mem_183_2_W0_mask)
  );
  split_mem_0_ext mem_183_3 (
    .R0_addr(mem_183_3_R0_addr),
    .R0_clk(mem_183_3_R0_clk),
    .R0_data(mem_183_3_R0_data),
    .R0_en(mem_183_3_R0_en),
    .W0_addr(mem_183_3_W0_addr),
    .W0_clk(mem_183_3_W0_clk),
    .W0_data(mem_183_3_W0_data),
    .W0_en(mem_183_3_W0_en),
    .W0_mask(mem_183_3_W0_mask)
  );
  split_mem_0_ext mem_183_4 (
    .R0_addr(mem_183_4_R0_addr),
    .R0_clk(mem_183_4_R0_clk),
    .R0_data(mem_183_4_R0_data),
    .R0_en(mem_183_4_R0_en),
    .W0_addr(mem_183_4_W0_addr),
    .W0_clk(mem_183_4_W0_clk),
    .W0_data(mem_183_4_W0_data),
    .W0_en(mem_183_4_W0_en),
    .W0_mask(mem_183_4_W0_mask)
  );
  split_mem_0_ext mem_183_5 (
    .R0_addr(mem_183_5_R0_addr),
    .R0_clk(mem_183_5_R0_clk),
    .R0_data(mem_183_5_R0_data),
    .R0_en(mem_183_5_R0_en),
    .W0_addr(mem_183_5_W0_addr),
    .W0_clk(mem_183_5_W0_clk),
    .W0_data(mem_183_5_W0_data),
    .W0_en(mem_183_5_W0_en),
    .W0_mask(mem_183_5_W0_mask)
  );
  split_mem_0_ext mem_183_6 (
    .R0_addr(mem_183_6_R0_addr),
    .R0_clk(mem_183_6_R0_clk),
    .R0_data(mem_183_6_R0_data),
    .R0_en(mem_183_6_R0_en),
    .W0_addr(mem_183_6_W0_addr),
    .W0_clk(mem_183_6_W0_clk),
    .W0_data(mem_183_6_W0_data),
    .W0_en(mem_183_6_W0_en),
    .W0_mask(mem_183_6_W0_mask)
  );
  split_mem_0_ext mem_183_7 (
    .R0_addr(mem_183_7_R0_addr),
    .R0_clk(mem_183_7_R0_clk),
    .R0_data(mem_183_7_R0_data),
    .R0_en(mem_183_7_R0_en),
    .W0_addr(mem_183_7_W0_addr),
    .W0_clk(mem_183_7_W0_clk),
    .W0_data(mem_183_7_W0_data),
    .W0_en(mem_183_7_W0_en),
    .W0_mask(mem_183_7_W0_mask)
  );
  split_mem_0_ext mem_184_0 (
    .R0_addr(mem_184_0_R0_addr),
    .R0_clk(mem_184_0_R0_clk),
    .R0_data(mem_184_0_R0_data),
    .R0_en(mem_184_0_R0_en),
    .W0_addr(mem_184_0_W0_addr),
    .W0_clk(mem_184_0_W0_clk),
    .W0_data(mem_184_0_W0_data),
    .W0_en(mem_184_0_W0_en),
    .W0_mask(mem_184_0_W0_mask)
  );
  split_mem_0_ext mem_184_1 (
    .R0_addr(mem_184_1_R0_addr),
    .R0_clk(mem_184_1_R0_clk),
    .R0_data(mem_184_1_R0_data),
    .R0_en(mem_184_1_R0_en),
    .W0_addr(mem_184_1_W0_addr),
    .W0_clk(mem_184_1_W0_clk),
    .W0_data(mem_184_1_W0_data),
    .W0_en(mem_184_1_W0_en),
    .W0_mask(mem_184_1_W0_mask)
  );
  split_mem_0_ext mem_184_2 (
    .R0_addr(mem_184_2_R0_addr),
    .R0_clk(mem_184_2_R0_clk),
    .R0_data(mem_184_2_R0_data),
    .R0_en(mem_184_2_R0_en),
    .W0_addr(mem_184_2_W0_addr),
    .W0_clk(mem_184_2_W0_clk),
    .W0_data(mem_184_2_W0_data),
    .W0_en(mem_184_2_W0_en),
    .W0_mask(mem_184_2_W0_mask)
  );
  split_mem_0_ext mem_184_3 (
    .R0_addr(mem_184_3_R0_addr),
    .R0_clk(mem_184_3_R0_clk),
    .R0_data(mem_184_3_R0_data),
    .R0_en(mem_184_3_R0_en),
    .W0_addr(mem_184_3_W0_addr),
    .W0_clk(mem_184_3_W0_clk),
    .W0_data(mem_184_3_W0_data),
    .W0_en(mem_184_3_W0_en),
    .W0_mask(mem_184_3_W0_mask)
  );
  split_mem_0_ext mem_184_4 (
    .R0_addr(mem_184_4_R0_addr),
    .R0_clk(mem_184_4_R0_clk),
    .R0_data(mem_184_4_R0_data),
    .R0_en(mem_184_4_R0_en),
    .W0_addr(mem_184_4_W0_addr),
    .W0_clk(mem_184_4_W0_clk),
    .W0_data(mem_184_4_W0_data),
    .W0_en(mem_184_4_W0_en),
    .W0_mask(mem_184_4_W0_mask)
  );
  split_mem_0_ext mem_184_5 (
    .R0_addr(mem_184_5_R0_addr),
    .R0_clk(mem_184_5_R0_clk),
    .R0_data(mem_184_5_R0_data),
    .R0_en(mem_184_5_R0_en),
    .W0_addr(mem_184_5_W0_addr),
    .W0_clk(mem_184_5_W0_clk),
    .W0_data(mem_184_5_W0_data),
    .W0_en(mem_184_5_W0_en),
    .W0_mask(mem_184_5_W0_mask)
  );
  split_mem_0_ext mem_184_6 (
    .R0_addr(mem_184_6_R0_addr),
    .R0_clk(mem_184_6_R0_clk),
    .R0_data(mem_184_6_R0_data),
    .R0_en(mem_184_6_R0_en),
    .W0_addr(mem_184_6_W0_addr),
    .W0_clk(mem_184_6_W0_clk),
    .W0_data(mem_184_6_W0_data),
    .W0_en(mem_184_6_W0_en),
    .W0_mask(mem_184_6_W0_mask)
  );
  split_mem_0_ext mem_184_7 (
    .R0_addr(mem_184_7_R0_addr),
    .R0_clk(mem_184_7_R0_clk),
    .R0_data(mem_184_7_R0_data),
    .R0_en(mem_184_7_R0_en),
    .W0_addr(mem_184_7_W0_addr),
    .W0_clk(mem_184_7_W0_clk),
    .W0_data(mem_184_7_W0_data),
    .W0_en(mem_184_7_W0_en),
    .W0_mask(mem_184_7_W0_mask)
  );
  split_mem_0_ext mem_185_0 (
    .R0_addr(mem_185_0_R0_addr),
    .R0_clk(mem_185_0_R0_clk),
    .R0_data(mem_185_0_R0_data),
    .R0_en(mem_185_0_R0_en),
    .W0_addr(mem_185_0_W0_addr),
    .W0_clk(mem_185_0_W0_clk),
    .W0_data(mem_185_0_W0_data),
    .W0_en(mem_185_0_W0_en),
    .W0_mask(mem_185_0_W0_mask)
  );
  split_mem_0_ext mem_185_1 (
    .R0_addr(mem_185_1_R0_addr),
    .R0_clk(mem_185_1_R0_clk),
    .R0_data(mem_185_1_R0_data),
    .R0_en(mem_185_1_R0_en),
    .W0_addr(mem_185_1_W0_addr),
    .W0_clk(mem_185_1_W0_clk),
    .W0_data(mem_185_1_W0_data),
    .W0_en(mem_185_1_W0_en),
    .W0_mask(mem_185_1_W0_mask)
  );
  split_mem_0_ext mem_185_2 (
    .R0_addr(mem_185_2_R0_addr),
    .R0_clk(mem_185_2_R0_clk),
    .R0_data(mem_185_2_R0_data),
    .R0_en(mem_185_2_R0_en),
    .W0_addr(mem_185_2_W0_addr),
    .W0_clk(mem_185_2_W0_clk),
    .W0_data(mem_185_2_W0_data),
    .W0_en(mem_185_2_W0_en),
    .W0_mask(mem_185_2_W0_mask)
  );
  split_mem_0_ext mem_185_3 (
    .R0_addr(mem_185_3_R0_addr),
    .R0_clk(mem_185_3_R0_clk),
    .R0_data(mem_185_3_R0_data),
    .R0_en(mem_185_3_R0_en),
    .W0_addr(mem_185_3_W0_addr),
    .W0_clk(mem_185_3_W0_clk),
    .W0_data(mem_185_3_W0_data),
    .W0_en(mem_185_3_W0_en),
    .W0_mask(mem_185_3_W0_mask)
  );
  split_mem_0_ext mem_185_4 (
    .R0_addr(mem_185_4_R0_addr),
    .R0_clk(mem_185_4_R0_clk),
    .R0_data(mem_185_4_R0_data),
    .R0_en(mem_185_4_R0_en),
    .W0_addr(mem_185_4_W0_addr),
    .W0_clk(mem_185_4_W0_clk),
    .W0_data(mem_185_4_W0_data),
    .W0_en(mem_185_4_W0_en),
    .W0_mask(mem_185_4_W0_mask)
  );
  split_mem_0_ext mem_185_5 (
    .R0_addr(mem_185_5_R0_addr),
    .R0_clk(mem_185_5_R0_clk),
    .R0_data(mem_185_5_R0_data),
    .R0_en(mem_185_5_R0_en),
    .W0_addr(mem_185_5_W0_addr),
    .W0_clk(mem_185_5_W0_clk),
    .W0_data(mem_185_5_W0_data),
    .W0_en(mem_185_5_W0_en),
    .W0_mask(mem_185_5_W0_mask)
  );
  split_mem_0_ext mem_185_6 (
    .R0_addr(mem_185_6_R0_addr),
    .R0_clk(mem_185_6_R0_clk),
    .R0_data(mem_185_6_R0_data),
    .R0_en(mem_185_6_R0_en),
    .W0_addr(mem_185_6_W0_addr),
    .W0_clk(mem_185_6_W0_clk),
    .W0_data(mem_185_6_W0_data),
    .W0_en(mem_185_6_W0_en),
    .W0_mask(mem_185_6_W0_mask)
  );
  split_mem_0_ext mem_185_7 (
    .R0_addr(mem_185_7_R0_addr),
    .R0_clk(mem_185_7_R0_clk),
    .R0_data(mem_185_7_R0_data),
    .R0_en(mem_185_7_R0_en),
    .W0_addr(mem_185_7_W0_addr),
    .W0_clk(mem_185_7_W0_clk),
    .W0_data(mem_185_7_W0_data),
    .W0_en(mem_185_7_W0_en),
    .W0_mask(mem_185_7_W0_mask)
  );
  split_mem_0_ext mem_186_0 (
    .R0_addr(mem_186_0_R0_addr),
    .R0_clk(mem_186_0_R0_clk),
    .R0_data(mem_186_0_R0_data),
    .R0_en(mem_186_0_R0_en),
    .W0_addr(mem_186_0_W0_addr),
    .W0_clk(mem_186_0_W0_clk),
    .W0_data(mem_186_0_W0_data),
    .W0_en(mem_186_0_W0_en),
    .W0_mask(mem_186_0_W0_mask)
  );
  split_mem_0_ext mem_186_1 (
    .R0_addr(mem_186_1_R0_addr),
    .R0_clk(mem_186_1_R0_clk),
    .R0_data(mem_186_1_R0_data),
    .R0_en(mem_186_1_R0_en),
    .W0_addr(mem_186_1_W0_addr),
    .W0_clk(mem_186_1_W0_clk),
    .W0_data(mem_186_1_W0_data),
    .W0_en(mem_186_1_W0_en),
    .W0_mask(mem_186_1_W0_mask)
  );
  split_mem_0_ext mem_186_2 (
    .R0_addr(mem_186_2_R0_addr),
    .R0_clk(mem_186_2_R0_clk),
    .R0_data(mem_186_2_R0_data),
    .R0_en(mem_186_2_R0_en),
    .W0_addr(mem_186_2_W0_addr),
    .W0_clk(mem_186_2_W0_clk),
    .W0_data(mem_186_2_W0_data),
    .W0_en(mem_186_2_W0_en),
    .W0_mask(mem_186_2_W0_mask)
  );
  split_mem_0_ext mem_186_3 (
    .R0_addr(mem_186_3_R0_addr),
    .R0_clk(mem_186_3_R0_clk),
    .R0_data(mem_186_3_R0_data),
    .R0_en(mem_186_3_R0_en),
    .W0_addr(mem_186_3_W0_addr),
    .W0_clk(mem_186_3_W0_clk),
    .W0_data(mem_186_3_W0_data),
    .W0_en(mem_186_3_W0_en),
    .W0_mask(mem_186_3_W0_mask)
  );
  split_mem_0_ext mem_186_4 (
    .R0_addr(mem_186_4_R0_addr),
    .R0_clk(mem_186_4_R0_clk),
    .R0_data(mem_186_4_R0_data),
    .R0_en(mem_186_4_R0_en),
    .W0_addr(mem_186_4_W0_addr),
    .W0_clk(mem_186_4_W0_clk),
    .W0_data(mem_186_4_W0_data),
    .W0_en(mem_186_4_W0_en),
    .W0_mask(mem_186_4_W0_mask)
  );
  split_mem_0_ext mem_186_5 (
    .R0_addr(mem_186_5_R0_addr),
    .R0_clk(mem_186_5_R0_clk),
    .R0_data(mem_186_5_R0_data),
    .R0_en(mem_186_5_R0_en),
    .W0_addr(mem_186_5_W0_addr),
    .W0_clk(mem_186_5_W0_clk),
    .W0_data(mem_186_5_W0_data),
    .W0_en(mem_186_5_W0_en),
    .W0_mask(mem_186_5_W0_mask)
  );
  split_mem_0_ext mem_186_6 (
    .R0_addr(mem_186_6_R0_addr),
    .R0_clk(mem_186_6_R0_clk),
    .R0_data(mem_186_6_R0_data),
    .R0_en(mem_186_6_R0_en),
    .W0_addr(mem_186_6_W0_addr),
    .W0_clk(mem_186_6_W0_clk),
    .W0_data(mem_186_6_W0_data),
    .W0_en(mem_186_6_W0_en),
    .W0_mask(mem_186_6_W0_mask)
  );
  split_mem_0_ext mem_186_7 (
    .R0_addr(mem_186_7_R0_addr),
    .R0_clk(mem_186_7_R0_clk),
    .R0_data(mem_186_7_R0_data),
    .R0_en(mem_186_7_R0_en),
    .W0_addr(mem_186_7_W0_addr),
    .W0_clk(mem_186_7_W0_clk),
    .W0_data(mem_186_7_W0_data),
    .W0_en(mem_186_7_W0_en),
    .W0_mask(mem_186_7_W0_mask)
  );
  split_mem_0_ext mem_187_0 (
    .R0_addr(mem_187_0_R0_addr),
    .R0_clk(mem_187_0_R0_clk),
    .R0_data(mem_187_0_R0_data),
    .R0_en(mem_187_0_R0_en),
    .W0_addr(mem_187_0_W0_addr),
    .W0_clk(mem_187_0_W0_clk),
    .W0_data(mem_187_0_W0_data),
    .W0_en(mem_187_0_W0_en),
    .W0_mask(mem_187_0_W0_mask)
  );
  split_mem_0_ext mem_187_1 (
    .R0_addr(mem_187_1_R0_addr),
    .R0_clk(mem_187_1_R0_clk),
    .R0_data(mem_187_1_R0_data),
    .R0_en(mem_187_1_R0_en),
    .W0_addr(mem_187_1_W0_addr),
    .W0_clk(mem_187_1_W0_clk),
    .W0_data(mem_187_1_W0_data),
    .W0_en(mem_187_1_W0_en),
    .W0_mask(mem_187_1_W0_mask)
  );
  split_mem_0_ext mem_187_2 (
    .R0_addr(mem_187_2_R0_addr),
    .R0_clk(mem_187_2_R0_clk),
    .R0_data(mem_187_2_R0_data),
    .R0_en(mem_187_2_R0_en),
    .W0_addr(mem_187_2_W0_addr),
    .W0_clk(mem_187_2_W0_clk),
    .W0_data(mem_187_2_W0_data),
    .W0_en(mem_187_2_W0_en),
    .W0_mask(mem_187_2_W0_mask)
  );
  split_mem_0_ext mem_187_3 (
    .R0_addr(mem_187_3_R0_addr),
    .R0_clk(mem_187_3_R0_clk),
    .R0_data(mem_187_3_R0_data),
    .R0_en(mem_187_3_R0_en),
    .W0_addr(mem_187_3_W0_addr),
    .W0_clk(mem_187_3_W0_clk),
    .W0_data(mem_187_3_W0_data),
    .W0_en(mem_187_3_W0_en),
    .W0_mask(mem_187_3_W0_mask)
  );
  split_mem_0_ext mem_187_4 (
    .R0_addr(mem_187_4_R0_addr),
    .R0_clk(mem_187_4_R0_clk),
    .R0_data(mem_187_4_R0_data),
    .R0_en(mem_187_4_R0_en),
    .W0_addr(mem_187_4_W0_addr),
    .W0_clk(mem_187_4_W0_clk),
    .W0_data(mem_187_4_W0_data),
    .W0_en(mem_187_4_W0_en),
    .W0_mask(mem_187_4_W0_mask)
  );
  split_mem_0_ext mem_187_5 (
    .R0_addr(mem_187_5_R0_addr),
    .R0_clk(mem_187_5_R0_clk),
    .R0_data(mem_187_5_R0_data),
    .R0_en(mem_187_5_R0_en),
    .W0_addr(mem_187_5_W0_addr),
    .W0_clk(mem_187_5_W0_clk),
    .W0_data(mem_187_5_W0_data),
    .W0_en(mem_187_5_W0_en),
    .W0_mask(mem_187_5_W0_mask)
  );
  split_mem_0_ext mem_187_6 (
    .R0_addr(mem_187_6_R0_addr),
    .R0_clk(mem_187_6_R0_clk),
    .R0_data(mem_187_6_R0_data),
    .R0_en(mem_187_6_R0_en),
    .W0_addr(mem_187_6_W0_addr),
    .W0_clk(mem_187_6_W0_clk),
    .W0_data(mem_187_6_W0_data),
    .W0_en(mem_187_6_W0_en),
    .W0_mask(mem_187_6_W0_mask)
  );
  split_mem_0_ext mem_187_7 (
    .R0_addr(mem_187_7_R0_addr),
    .R0_clk(mem_187_7_R0_clk),
    .R0_data(mem_187_7_R0_data),
    .R0_en(mem_187_7_R0_en),
    .W0_addr(mem_187_7_W0_addr),
    .W0_clk(mem_187_7_W0_clk),
    .W0_data(mem_187_7_W0_data),
    .W0_en(mem_187_7_W0_en),
    .W0_mask(mem_187_7_W0_mask)
  );
  split_mem_0_ext mem_188_0 (
    .R0_addr(mem_188_0_R0_addr),
    .R0_clk(mem_188_0_R0_clk),
    .R0_data(mem_188_0_R0_data),
    .R0_en(mem_188_0_R0_en),
    .W0_addr(mem_188_0_W0_addr),
    .W0_clk(mem_188_0_W0_clk),
    .W0_data(mem_188_0_W0_data),
    .W0_en(mem_188_0_W0_en),
    .W0_mask(mem_188_0_W0_mask)
  );
  split_mem_0_ext mem_188_1 (
    .R0_addr(mem_188_1_R0_addr),
    .R0_clk(mem_188_1_R0_clk),
    .R0_data(mem_188_1_R0_data),
    .R0_en(mem_188_1_R0_en),
    .W0_addr(mem_188_1_W0_addr),
    .W0_clk(mem_188_1_W0_clk),
    .W0_data(mem_188_1_W0_data),
    .W0_en(mem_188_1_W0_en),
    .W0_mask(mem_188_1_W0_mask)
  );
  split_mem_0_ext mem_188_2 (
    .R0_addr(mem_188_2_R0_addr),
    .R0_clk(mem_188_2_R0_clk),
    .R0_data(mem_188_2_R0_data),
    .R0_en(mem_188_2_R0_en),
    .W0_addr(mem_188_2_W0_addr),
    .W0_clk(mem_188_2_W0_clk),
    .W0_data(mem_188_2_W0_data),
    .W0_en(mem_188_2_W0_en),
    .W0_mask(mem_188_2_W0_mask)
  );
  split_mem_0_ext mem_188_3 (
    .R0_addr(mem_188_3_R0_addr),
    .R0_clk(mem_188_3_R0_clk),
    .R0_data(mem_188_3_R0_data),
    .R0_en(mem_188_3_R0_en),
    .W0_addr(mem_188_3_W0_addr),
    .W0_clk(mem_188_3_W0_clk),
    .W0_data(mem_188_3_W0_data),
    .W0_en(mem_188_3_W0_en),
    .W0_mask(mem_188_3_W0_mask)
  );
  split_mem_0_ext mem_188_4 (
    .R0_addr(mem_188_4_R0_addr),
    .R0_clk(mem_188_4_R0_clk),
    .R0_data(mem_188_4_R0_data),
    .R0_en(mem_188_4_R0_en),
    .W0_addr(mem_188_4_W0_addr),
    .W0_clk(mem_188_4_W0_clk),
    .W0_data(mem_188_4_W0_data),
    .W0_en(mem_188_4_W0_en),
    .W0_mask(mem_188_4_W0_mask)
  );
  split_mem_0_ext mem_188_5 (
    .R0_addr(mem_188_5_R0_addr),
    .R0_clk(mem_188_5_R0_clk),
    .R0_data(mem_188_5_R0_data),
    .R0_en(mem_188_5_R0_en),
    .W0_addr(mem_188_5_W0_addr),
    .W0_clk(mem_188_5_W0_clk),
    .W0_data(mem_188_5_W0_data),
    .W0_en(mem_188_5_W0_en),
    .W0_mask(mem_188_5_W0_mask)
  );
  split_mem_0_ext mem_188_6 (
    .R0_addr(mem_188_6_R0_addr),
    .R0_clk(mem_188_6_R0_clk),
    .R0_data(mem_188_6_R0_data),
    .R0_en(mem_188_6_R0_en),
    .W0_addr(mem_188_6_W0_addr),
    .W0_clk(mem_188_6_W0_clk),
    .W0_data(mem_188_6_W0_data),
    .W0_en(mem_188_6_W0_en),
    .W0_mask(mem_188_6_W0_mask)
  );
  split_mem_0_ext mem_188_7 (
    .R0_addr(mem_188_7_R0_addr),
    .R0_clk(mem_188_7_R0_clk),
    .R0_data(mem_188_7_R0_data),
    .R0_en(mem_188_7_R0_en),
    .W0_addr(mem_188_7_W0_addr),
    .W0_clk(mem_188_7_W0_clk),
    .W0_data(mem_188_7_W0_data),
    .W0_en(mem_188_7_W0_en),
    .W0_mask(mem_188_7_W0_mask)
  );
  split_mem_0_ext mem_189_0 (
    .R0_addr(mem_189_0_R0_addr),
    .R0_clk(mem_189_0_R0_clk),
    .R0_data(mem_189_0_R0_data),
    .R0_en(mem_189_0_R0_en),
    .W0_addr(mem_189_0_W0_addr),
    .W0_clk(mem_189_0_W0_clk),
    .W0_data(mem_189_0_W0_data),
    .W0_en(mem_189_0_W0_en),
    .W0_mask(mem_189_0_W0_mask)
  );
  split_mem_0_ext mem_189_1 (
    .R0_addr(mem_189_1_R0_addr),
    .R0_clk(mem_189_1_R0_clk),
    .R0_data(mem_189_1_R0_data),
    .R0_en(mem_189_1_R0_en),
    .W0_addr(mem_189_1_W0_addr),
    .W0_clk(mem_189_1_W0_clk),
    .W0_data(mem_189_1_W0_data),
    .W0_en(mem_189_1_W0_en),
    .W0_mask(mem_189_1_W0_mask)
  );
  split_mem_0_ext mem_189_2 (
    .R0_addr(mem_189_2_R0_addr),
    .R0_clk(mem_189_2_R0_clk),
    .R0_data(mem_189_2_R0_data),
    .R0_en(mem_189_2_R0_en),
    .W0_addr(mem_189_2_W0_addr),
    .W0_clk(mem_189_2_W0_clk),
    .W0_data(mem_189_2_W0_data),
    .W0_en(mem_189_2_W0_en),
    .W0_mask(mem_189_2_W0_mask)
  );
  split_mem_0_ext mem_189_3 (
    .R0_addr(mem_189_3_R0_addr),
    .R0_clk(mem_189_3_R0_clk),
    .R0_data(mem_189_3_R0_data),
    .R0_en(mem_189_3_R0_en),
    .W0_addr(mem_189_3_W0_addr),
    .W0_clk(mem_189_3_W0_clk),
    .W0_data(mem_189_3_W0_data),
    .W0_en(mem_189_3_W0_en),
    .W0_mask(mem_189_3_W0_mask)
  );
  split_mem_0_ext mem_189_4 (
    .R0_addr(mem_189_4_R0_addr),
    .R0_clk(mem_189_4_R0_clk),
    .R0_data(mem_189_4_R0_data),
    .R0_en(mem_189_4_R0_en),
    .W0_addr(mem_189_4_W0_addr),
    .W0_clk(mem_189_4_W0_clk),
    .W0_data(mem_189_4_W0_data),
    .W0_en(mem_189_4_W0_en),
    .W0_mask(mem_189_4_W0_mask)
  );
  split_mem_0_ext mem_189_5 (
    .R0_addr(mem_189_5_R0_addr),
    .R0_clk(mem_189_5_R0_clk),
    .R0_data(mem_189_5_R0_data),
    .R0_en(mem_189_5_R0_en),
    .W0_addr(mem_189_5_W0_addr),
    .W0_clk(mem_189_5_W0_clk),
    .W0_data(mem_189_5_W0_data),
    .W0_en(mem_189_5_W0_en),
    .W0_mask(mem_189_5_W0_mask)
  );
  split_mem_0_ext mem_189_6 (
    .R0_addr(mem_189_6_R0_addr),
    .R0_clk(mem_189_6_R0_clk),
    .R0_data(mem_189_6_R0_data),
    .R0_en(mem_189_6_R0_en),
    .W0_addr(mem_189_6_W0_addr),
    .W0_clk(mem_189_6_W0_clk),
    .W0_data(mem_189_6_W0_data),
    .W0_en(mem_189_6_W0_en),
    .W0_mask(mem_189_6_W0_mask)
  );
  split_mem_0_ext mem_189_7 (
    .R0_addr(mem_189_7_R0_addr),
    .R0_clk(mem_189_7_R0_clk),
    .R0_data(mem_189_7_R0_data),
    .R0_en(mem_189_7_R0_en),
    .W0_addr(mem_189_7_W0_addr),
    .W0_clk(mem_189_7_W0_clk),
    .W0_data(mem_189_7_W0_data),
    .W0_en(mem_189_7_W0_en),
    .W0_mask(mem_189_7_W0_mask)
  );
  split_mem_0_ext mem_190_0 (
    .R0_addr(mem_190_0_R0_addr),
    .R0_clk(mem_190_0_R0_clk),
    .R0_data(mem_190_0_R0_data),
    .R0_en(mem_190_0_R0_en),
    .W0_addr(mem_190_0_W0_addr),
    .W0_clk(mem_190_0_W0_clk),
    .W0_data(mem_190_0_W0_data),
    .W0_en(mem_190_0_W0_en),
    .W0_mask(mem_190_0_W0_mask)
  );
  split_mem_0_ext mem_190_1 (
    .R0_addr(mem_190_1_R0_addr),
    .R0_clk(mem_190_1_R0_clk),
    .R0_data(mem_190_1_R0_data),
    .R0_en(mem_190_1_R0_en),
    .W0_addr(mem_190_1_W0_addr),
    .W0_clk(mem_190_1_W0_clk),
    .W0_data(mem_190_1_W0_data),
    .W0_en(mem_190_1_W0_en),
    .W0_mask(mem_190_1_W0_mask)
  );
  split_mem_0_ext mem_190_2 (
    .R0_addr(mem_190_2_R0_addr),
    .R0_clk(mem_190_2_R0_clk),
    .R0_data(mem_190_2_R0_data),
    .R0_en(mem_190_2_R0_en),
    .W0_addr(mem_190_2_W0_addr),
    .W0_clk(mem_190_2_W0_clk),
    .W0_data(mem_190_2_W0_data),
    .W0_en(mem_190_2_W0_en),
    .W0_mask(mem_190_2_W0_mask)
  );
  split_mem_0_ext mem_190_3 (
    .R0_addr(mem_190_3_R0_addr),
    .R0_clk(mem_190_3_R0_clk),
    .R0_data(mem_190_3_R0_data),
    .R0_en(mem_190_3_R0_en),
    .W0_addr(mem_190_3_W0_addr),
    .W0_clk(mem_190_3_W0_clk),
    .W0_data(mem_190_3_W0_data),
    .W0_en(mem_190_3_W0_en),
    .W0_mask(mem_190_3_W0_mask)
  );
  split_mem_0_ext mem_190_4 (
    .R0_addr(mem_190_4_R0_addr),
    .R0_clk(mem_190_4_R0_clk),
    .R0_data(mem_190_4_R0_data),
    .R0_en(mem_190_4_R0_en),
    .W0_addr(mem_190_4_W0_addr),
    .W0_clk(mem_190_4_W0_clk),
    .W0_data(mem_190_4_W0_data),
    .W0_en(mem_190_4_W0_en),
    .W0_mask(mem_190_4_W0_mask)
  );
  split_mem_0_ext mem_190_5 (
    .R0_addr(mem_190_5_R0_addr),
    .R0_clk(mem_190_5_R0_clk),
    .R0_data(mem_190_5_R0_data),
    .R0_en(mem_190_5_R0_en),
    .W0_addr(mem_190_5_W0_addr),
    .W0_clk(mem_190_5_W0_clk),
    .W0_data(mem_190_5_W0_data),
    .W0_en(mem_190_5_W0_en),
    .W0_mask(mem_190_5_W0_mask)
  );
  split_mem_0_ext mem_190_6 (
    .R0_addr(mem_190_6_R0_addr),
    .R0_clk(mem_190_6_R0_clk),
    .R0_data(mem_190_6_R0_data),
    .R0_en(mem_190_6_R0_en),
    .W0_addr(mem_190_6_W0_addr),
    .W0_clk(mem_190_6_W0_clk),
    .W0_data(mem_190_6_W0_data),
    .W0_en(mem_190_6_W0_en),
    .W0_mask(mem_190_6_W0_mask)
  );
  split_mem_0_ext mem_190_7 (
    .R0_addr(mem_190_7_R0_addr),
    .R0_clk(mem_190_7_R0_clk),
    .R0_data(mem_190_7_R0_data),
    .R0_en(mem_190_7_R0_en),
    .W0_addr(mem_190_7_W0_addr),
    .W0_clk(mem_190_7_W0_clk),
    .W0_data(mem_190_7_W0_data),
    .W0_en(mem_190_7_W0_en),
    .W0_mask(mem_190_7_W0_mask)
  );
  split_mem_0_ext mem_191_0 (
    .R0_addr(mem_191_0_R0_addr),
    .R0_clk(mem_191_0_R0_clk),
    .R0_data(mem_191_0_R0_data),
    .R0_en(mem_191_0_R0_en),
    .W0_addr(mem_191_0_W0_addr),
    .W0_clk(mem_191_0_W0_clk),
    .W0_data(mem_191_0_W0_data),
    .W0_en(mem_191_0_W0_en),
    .W0_mask(mem_191_0_W0_mask)
  );
  split_mem_0_ext mem_191_1 (
    .R0_addr(mem_191_1_R0_addr),
    .R0_clk(mem_191_1_R0_clk),
    .R0_data(mem_191_1_R0_data),
    .R0_en(mem_191_1_R0_en),
    .W0_addr(mem_191_1_W0_addr),
    .W0_clk(mem_191_1_W0_clk),
    .W0_data(mem_191_1_W0_data),
    .W0_en(mem_191_1_W0_en),
    .W0_mask(mem_191_1_W0_mask)
  );
  split_mem_0_ext mem_191_2 (
    .R0_addr(mem_191_2_R0_addr),
    .R0_clk(mem_191_2_R0_clk),
    .R0_data(mem_191_2_R0_data),
    .R0_en(mem_191_2_R0_en),
    .W0_addr(mem_191_2_W0_addr),
    .W0_clk(mem_191_2_W0_clk),
    .W0_data(mem_191_2_W0_data),
    .W0_en(mem_191_2_W0_en),
    .W0_mask(mem_191_2_W0_mask)
  );
  split_mem_0_ext mem_191_3 (
    .R0_addr(mem_191_3_R0_addr),
    .R0_clk(mem_191_3_R0_clk),
    .R0_data(mem_191_3_R0_data),
    .R0_en(mem_191_3_R0_en),
    .W0_addr(mem_191_3_W0_addr),
    .W0_clk(mem_191_3_W0_clk),
    .W0_data(mem_191_3_W0_data),
    .W0_en(mem_191_3_W0_en),
    .W0_mask(mem_191_3_W0_mask)
  );
  split_mem_0_ext mem_191_4 (
    .R0_addr(mem_191_4_R0_addr),
    .R0_clk(mem_191_4_R0_clk),
    .R0_data(mem_191_4_R0_data),
    .R0_en(mem_191_4_R0_en),
    .W0_addr(mem_191_4_W0_addr),
    .W0_clk(mem_191_4_W0_clk),
    .W0_data(mem_191_4_W0_data),
    .W0_en(mem_191_4_W0_en),
    .W0_mask(mem_191_4_W0_mask)
  );
  split_mem_0_ext mem_191_5 (
    .R0_addr(mem_191_5_R0_addr),
    .R0_clk(mem_191_5_R0_clk),
    .R0_data(mem_191_5_R0_data),
    .R0_en(mem_191_5_R0_en),
    .W0_addr(mem_191_5_W0_addr),
    .W0_clk(mem_191_5_W0_clk),
    .W0_data(mem_191_5_W0_data),
    .W0_en(mem_191_5_W0_en),
    .W0_mask(mem_191_5_W0_mask)
  );
  split_mem_0_ext mem_191_6 (
    .R0_addr(mem_191_6_R0_addr),
    .R0_clk(mem_191_6_R0_clk),
    .R0_data(mem_191_6_R0_data),
    .R0_en(mem_191_6_R0_en),
    .W0_addr(mem_191_6_W0_addr),
    .W0_clk(mem_191_6_W0_clk),
    .W0_data(mem_191_6_W0_data),
    .W0_en(mem_191_6_W0_en),
    .W0_mask(mem_191_6_W0_mask)
  );
  split_mem_0_ext mem_191_7 (
    .R0_addr(mem_191_7_R0_addr),
    .R0_clk(mem_191_7_R0_clk),
    .R0_data(mem_191_7_R0_data),
    .R0_en(mem_191_7_R0_en),
    .W0_addr(mem_191_7_W0_addr),
    .W0_clk(mem_191_7_W0_clk),
    .W0_data(mem_191_7_W0_data),
    .W0_en(mem_191_7_W0_en),
    .W0_mask(mem_191_7_W0_mask)
  );
  split_mem_0_ext mem_192_0 (
    .R0_addr(mem_192_0_R0_addr),
    .R0_clk(mem_192_0_R0_clk),
    .R0_data(mem_192_0_R0_data),
    .R0_en(mem_192_0_R0_en),
    .W0_addr(mem_192_0_W0_addr),
    .W0_clk(mem_192_0_W0_clk),
    .W0_data(mem_192_0_W0_data),
    .W0_en(mem_192_0_W0_en),
    .W0_mask(mem_192_0_W0_mask)
  );
  split_mem_0_ext mem_192_1 (
    .R0_addr(mem_192_1_R0_addr),
    .R0_clk(mem_192_1_R0_clk),
    .R0_data(mem_192_1_R0_data),
    .R0_en(mem_192_1_R0_en),
    .W0_addr(mem_192_1_W0_addr),
    .W0_clk(mem_192_1_W0_clk),
    .W0_data(mem_192_1_W0_data),
    .W0_en(mem_192_1_W0_en),
    .W0_mask(mem_192_1_W0_mask)
  );
  split_mem_0_ext mem_192_2 (
    .R0_addr(mem_192_2_R0_addr),
    .R0_clk(mem_192_2_R0_clk),
    .R0_data(mem_192_2_R0_data),
    .R0_en(mem_192_2_R0_en),
    .W0_addr(mem_192_2_W0_addr),
    .W0_clk(mem_192_2_W0_clk),
    .W0_data(mem_192_2_W0_data),
    .W0_en(mem_192_2_W0_en),
    .W0_mask(mem_192_2_W0_mask)
  );
  split_mem_0_ext mem_192_3 (
    .R0_addr(mem_192_3_R0_addr),
    .R0_clk(mem_192_3_R0_clk),
    .R0_data(mem_192_3_R0_data),
    .R0_en(mem_192_3_R0_en),
    .W0_addr(mem_192_3_W0_addr),
    .W0_clk(mem_192_3_W0_clk),
    .W0_data(mem_192_3_W0_data),
    .W0_en(mem_192_3_W0_en),
    .W0_mask(mem_192_3_W0_mask)
  );
  split_mem_0_ext mem_192_4 (
    .R0_addr(mem_192_4_R0_addr),
    .R0_clk(mem_192_4_R0_clk),
    .R0_data(mem_192_4_R0_data),
    .R0_en(mem_192_4_R0_en),
    .W0_addr(mem_192_4_W0_addr),
    .W0_clk(mem_192_4_W0_clk),
    .W0_data(mem_192_4_W0_data),
    .W0_en(mem_192_4_W0_en),
    .W0_mask(mem_192_4_W0_mask)
  );
  split_mem_0_ext mem_192_5 (
    .R0_addr(mem_192_5_R0_addr),
    .R0_clk(mem_192_5_R0_clk),
    .R0_data(mem_192_5_R0_data),
    .R0_en(mem_192_5_R0_en),
    .W0_addr(mem_192_5_W0_addr),
    .W0_clk(mem_192_5_W0_clk),
    .W0_data(mem_192_5_W0_data),
    .W0_en(mem_192_5_W0_en),
    .W0_mask(mem_192_5_W0_mask)
  );
  split_mem_0_ext mem_192_6 (
    .R0_addr(mem_192_6_R0_addr),
    .R0_clk(mem_192_6_R0_clk),
    .R0_data(mem_192_6_R0_data),
    .R0_en(mem_192_6_R0_en),
    .W0_addr(mem_192_6_W0_addr),
    .W0_clk(mem_192_6_W0_clk),
    .W0_data(mem_192_6_W0_data),
    .W0_en(mem_192_6_W0_en),
    .W0_mask(mem_192_6_W0_mask)
  );
  split_mem_0_ext mem_192_7 (
    .R0_addr(mem_192_7_R0_addr),
    .R0_clk(mem_192_7_R0_clk),
    .R0_data(mem_192_7_R0_data),
    .R0_en(mem_192_7_R0_en),
    .W0_addr(mem_192_7_W0_addr),
    .W0_clk(mem_192_7_W0_clk),
    .W0_data(mem_192_7_W0_data),
    .W0_en(mem_192_7_W0_en),
    .W0_mask(mem_192_7_W0_mask)
  );
  split_mem_0_ext mem_193_0 (
    .R0_addr(mem_193_0_R0_addr),
    .R0_clk(mem_193_0_R0_clk),
    .R0_data(mem_193_0_R0_data),
    .R0_en(mem_193_0_R0_en),
    .W0_addr(mem_193_0_W0_addr),
    .W0_clk(mem_193_0_W0_clk),
    .W0_data(mem_193_0_W0_data),
    .W0_en(mem_193_0_W0_en),
    .W0_mask(mem_193_0_W0_mask)
  );
  split_mem_0_ext mem_193_1 (
    .R0_addr(mem_193_1_R0_addr),
    .R0_clk(mem_193_1_R0_clk),
    .R0_data(mem_193_1_R0_data),
    .R0_en(mem_193_1_R0_en),
    .W0_addr(mem_193_1_W0_addr),
    .W0_clk(mem_193_1_W0_clk),
    .W0_data(mem_193_1_W0_data),
    .W0_en(mem_193_1_W0_en),
    .W0_mask(mem_193_1_W0_mask)
  );
  split_mem_0_ext mem_193_2 (
    .R0_addr(mem_193_2_R0_addr),
    .R0_clk(mem_193_2_R0_clk),
    .R0_data(mem_193_2_R0_data),
    .R0_en(mem_193_2_R0_en),
    .W0_addr(mem_193_2_W0_addr),
    .W0_clk(mem_193_2_W0_clk),
    .W0_data(mem_193_2_W0_data),
    .W0_en(mem_193_2_W0_en),
    .W0_mask(mem_193_2_W0_mask)
  );
  split_mem_0_ext mem_193_3 (
    .R0_addr(mem_193_3_R0_addr),
    .R0_clk(mem_193_3_R0_clk),
    .R0_data(mem_193_3_R0_data),
    .R0_en(mem_193_3_R0_en),
    .W0_addr(mem_193_3_W0_addr),
    .W0_clk(mem_193_3_W0_clk),
    .W0_data(mem_193_3_W0_data),
    .W0_en(mem_193_3_W0_en),
    .W0_mask(mem_193_3_W0_mask)
  );
  split_mem_0_ext mem_193_4 (
    .R0_addr(mem_193_4_R0_addr),
    .R0_clk(mem_193_4_R0_clk),
    .R0_data(mem_193_4_R0_data),
    .R0_en(mem_193_4_R0_en),
    .W0_addr(mem_193_4_W0_addr),
    .W0_clk(mem_193_4_W0_clk),
    .W0_data(mem_193_4_W0_data),
    .W0_en(mem_193_4_W0_en),
    .W0_mask(mem_193_4_W0_mask)
  );
  split_mem_0_ext mem_193_5 (
    .R0_addr(mem_193_5_R0_addr),
    .R0_clk(mem_193_5_R0_clk),
    .R0_data(mem_193_5_R0_data),
    .R0_en(mem_193_5_R0_en),
    .W0_addr(mem_193_5_W0_addr),
    .W0_clk(mem_193_5_W0_clk),
    .W0_data(mem_193_5_W0_data),
    .W0_en(mem_193_5_W0_en),
    .W0_mask(mem_193_5_W0_mask)
  );
  split_mem_0_ext mem_193_6 (
    .R0_addr(mem_193_6_R0_addr),
    .R0_clk(mem_193_6_R0_clk),
    .R0_data(mem_193_6_R0_data),
    .R0_en(mem_193_6_R0_en),
    .W0_addr(mem_193_6_W0_addr),
    .W0_clk(mem_193_6_W0_clk),
    .W0_data(mem_193_6_W0_data),
    .W0_en(mem_193_6_W0_en),
    .W0_mask(mem_193_6_W0_mask)
  );
  split_mem_0_ext mem_193_7 (
    .R0_addr(mem_193_7_R0_addr),
    .R0_clk(mem_193_7_R0_clk),
    .R0_data(mem_193_7_R0_data),
    .R0_en(mem_193_7_R0_en),
    .W0_addr(mem_193_7_W0_addr),
    .W0_clk(mem_193_7_W0_clk),
    .W0_data(mem_193_7_W0_data),
    .W0_en(mem_193_7_W0_en),
    .W0_mask(mem_193_7_W0_mask)
  );
  split_mem_0_ext mem_194_0 (
    .R0_addr(mem_194_0_R0_addr),
    .R0_clk(mem_194_0_R0_clk),
    .R0_data(mem_194_0_R0_data),
    .R0_en(mem_194_0_R0_en),
    .W0_addr(mem_194_0_W0_addr),
    .W0_clk(mem_194_0_W0_clk),
    .W0_data(mem_194_0_W0_data),
    .W0_en(mem_194_0_W0_en),
    .W0_mask(mem_194_0_W0_mask)
  );
  split_mem_0_ext mem_194_1 (
    .R0_addr(mem_194_1_R0_addr),
    .R0_clk(mem_194_1_R0_clk),
    .R0_data(mem_194_1_R0_data),
    .R0_en(mem_194_1_R0_en),
    .W0_addr(mem_194_1_W0_addr),
    .W0_clk(mem_194_1_W0_clk),
    .W0_data(mem_194_1_W0_data),
    .W0_en(mem_194_1_W0_en),
    .W0_mask(mem_194_1_W0_mask)
  );
  split_mem_0_ext mem_194_2 (
    .R0_addr(mem_194_2_R0_addr),
    .R0_clk(mem_194_2_R0_clk),
    .R0_data(mem_194_2_R0_data),
    .R0_en(mem_194_2_R0_en),
    .W0_addr(mem_194_2_W0_addr),
    .W0_clk(mem_194_2_W0_clk),
    .W0_data(mem_194_2_W0_data),
    .W0_en(mem_194_2_W0_en),
    .W0_mask(mem_194_2_W0_mask)
  );
  split_mem_0_ext mem_194_3 (
    .R0_addr(mem_194_3_R0_addr),
    .R0_clk(mem_194_3_R0_clk),
    .R0_data(mem_194_3_R0_data),
    .R0_en(mem_194_3_R0_en),
    .W0_addr(mem_194_3_W0_addr),
    .W0_clk(mem_194_3_W0_clk),
    .W0_data(mem_194_3_W0_data),
    .W0_en(mem_194_3_W0_en),
    .W0_mask(mem_194_3_W0_mask)
  );
  split_mem_0_ext mem_194_4 (
    .R0_addr(mem_194_4_R0_addr),
    .R0_clk(mem_194_4_R0_clk),
    .R0_data(mem_194_4_R0_data),
    .R0_en(mem_194_4_R0_en),
    .W0_addr(mem_194_4_W0_addr),
    .W0_clk(mem_194_4_W0_clk),
    .W0_data(mem_194_4_W0_data),
    .W0_en(mem_194_4_W0_en),
    .W0_mask(mem_194_4_W0_mask)
  );
  split_mem_0_ext mem_194_5 (
    .R0_addr(mem_194_5_R0_addr),
    .R0_clk(mem_194_5_R0_clk),
    .R0_data(mem_194_5_R0_data),
    .R0_en(mem_194_5_R0_en),
    .W0_addr(mem_194_5_W0_addr),
    .W0_clk(mem_194_5_W0_clk),
    .W0_data(mem_194_5_W0_data),
    .W0_en(mem_194_5_W0_en),
    .W0_mask(mem_194_5_W0_mask)
  );
  split_mem_0_ext mem_194_6 (
    .R0_addr(mem_194_6_R0_addr),
    .R0_clk(mem_194_6_R0_clk),
    .R0_data(mem_194_6_R0_data),
    .R0_en(mem_194_6_R0_en),
    .W0_addr(mem_194_6_W0_addr),
    .W0_clk(mem_194_6_W0_clk),
    .W0_data(mem_194_6_W0_data),
    .W0_en(mem_194_6_W0_en),
    .W0_mask(mem_194_6_W0_mask)
  );
  split_mem_0_ext mem_194_7 (
    .R0_addr(mem_194_7_R0_addr),
    .R0_clk(mem_194_7_R0_clk),
    .R0_data(mem_194_7_R0_data),
    .R0_en(mem_194_7_R0_en),
    .W0_addr(mem_194_7_W0_addr),
    .W0_clk(mem_194_7_W0_clk),
    .W0_data(mem_194_7_W0_data),
    .W0_en(mem_194_7_W0_en),
    .W0_mask(mem_194_7_W0_mask)
  );
  split_mem_0_ext mem_195_0 (
    .R0_addr(mem_195_0_R0_addr),
    .R0_clk(mem_195_0_R0_clk),
    .R0_data(mem_195_0_R0_data),
    .R0_en(mem_195_0_R0_en),
    .W0_addr(mem_195_0_W0_addr),
    .W0_clk(mem_195_0_W0_clk),
    .W0_data(mem_195_0_W0_data),
    .W0_en(mem_195_0_W0_en),
    .W0_mask(mem_195_0_W0_mask)
  );
  split_mem_0_ext mem_195_1 (
    .R0_addr(mem_195_1_R0_addr),
    .R0_clk(mem_195_1_R0_clk),
    .R0_data(mem_195_1_R0_data),
    .R0_en(mem_195_1_R0_en),
    .W0_addr(mem_195_1_W0_addr),
    .W0_clk(mem_195_1_W0_clk),
    .W0_data(mem_195_1_W0_data),
    .W0_en(mem_195_1_W0_en),
    .W0_mask(mem_195_1_W0_mask)
  );
  split_mem_0_ext mem_195_2 (
    .R0_addr(mem_195_2_R0_addr),
    .R0_clk(mem_195_2_R0_clk),
    .R0_data(mem_195_2_R0_data),
    .R0_en(mem_195_2_R0_en),
    .W0_addr(mem_195_2_W0_addr),
    .W0_clk(mem_195_2_W0_clk),
    .W0_data(mem_195_2_W0_data),
    .W0_en(mem_195_2_W0_en),
    .W0_mask(mem_195_2_W0_mask)
  );
  split_mem_0_ext mem_195_3 (
    .R0_addr(mem_195_3_R0_addr),
    .R0_clk(mem_195_3_R0_clk),
    .R0_data(mem_195_3_R0_data),
    .R0_en(mem_195_3_R0_en),
    .W0_addr(mem_195_3_W0_addr),
    .W0_clk(mem_195_3_W0_clk),
    .W0_data(mem_195_3_W0_data),
    .W0_en(mem_195_3_W0_en),
    .W0_mask(mem_195_3_W0_mask)
  );
  split_mem_0_ext mem_195_4 (
    .R0_addr(mem_195_4_R0_addr),
    .R0_clk(mem_195_4_R0_clk),
    .R0_data(mem_195_4_R0_data),
    .R0_en(mem_195_4_R0_en),
    .W0_addr(mem_195_4_W0_addr),
    .W0_clk(mem_195_4_W0_clk),
    .W0_data(mem_195_4_W0_data),
    .W0_en(mem_195_4_W0_en),
    .W0_mask(mem_195_4_W0_mask)
  );
  split_mem_0_ext mem_195_5 (
    .R0_addr(mem_195_5_R0_addr),
    .R0_clk(mem_195_5_R0_clk),
    .R0_data(mem_195_5_R0_data),
    .R0_en(mem_195_5_R0_en),
    .W0_addr(mem_195_5_W0_addr),
    .W0_clk(mem_195_5_W0_clk),
    .W0_data(mem_195_5_W0_data),
    .W0_en(mem_195_5_W0_en),
    .W0_mask(mem_195_5_W0_mask)
  );
  split_mem_0_ext mem_195_6 (
    .R0_addr(mem_195_6_R0_addr),
    .R0_clk(mem_195_6_R0_clk),
    .R0_data(mem_195_6_R0_data),
    .R0_en(mem_195_6_R0_en),
    .W0_addr(mem_195_6_W0_addr),
    .W0_clk(mem_195_6_W0_clk),
    .W0_data(mem_195_6_W0_data),
    .W0_en(mem_195_6_W0_en),
    .W0_mask(mem_195_6_W0_mask)
  );
  split_mem_0_ext mem_195_7 (
    .R0_addr(mem_195_7_R0_addr),
    .R0_clk(mem_195_7_R0_clk),
    .R0_data(mem_195_7_R0_data),
    .R0_en(mem_195_7_R0_en),
    .W0_addr(mem_195_7_W0_addr),
    .W0_clk(mem_195_7_W0_clk),
    .W0_data(mem_195_7_W0_data),
    .W0_en(mem_195_7_W0_en),
    .W0_mask(mem_195_7_W0_mask)
  );
  split_mem_0_ext mem_196_0 (
    .R0_addr(mem_196_0_R0_addr),
    .R0_clk(mem_196_0_R0_clk),
    .R0_data(mem_196_0_R0_data),
    .R0_en(mem_196_0_R0_en),
    .W0_addr(mem_196_0_W0_addr),
    .W0_clk(mem_196_0_W0_clk),
    .W0_data(mem_196_0_W0_data),
    .W0_en(mem_196_0_W0_en),
    .W0_mask(mem_196_0_W0_mask)
  );
  split_mem_0_ext mem_196_1 (
    .R0_addr(mem_196_1_R0_addr),
    .R0_clk(mem_196_1_R0_clk),
    .R0_data(mem_196_1_R0_data),
    .R0_en(mem_196_1_R0_en),
    .W0_addr(mem_196_1_W0_addr),
    .W0_clk(mem_196_1_W0_clk),
    .W0_data(mem_196_1_W0_data),
    .W0_en(mem_196_1_W0_en),
    .W0_mask(mem_196_1_W0_mask)
  );
  split_mem_0_ext mem_196_2 (
    .R0_addr(mem_196_2_R0_addr),
    .R0_clk(mem_196_2_R0_clk),
    .R0_data(mem_196_2_R0_data),
    .R0_en(mem_196_2_R0_en),
    .W0_addr(mem_196_2_W0_addr),
    .W0_clk(mem_196_2_W0_clk),
    .W0_data(mem_196_2_W0_data),
    .W0_en(mem_196_2_W0_en),
    .W0_mask(mem_196_2_W0_mask)
  );
  split_mem_0_ext mem_196_3 (
    .R0_addr(mem_196_3_R0_addr),
    .R0_clk(mem_196_3_R0_clk),
    .R0_data(mem_196_3_R0_data),
    .R0_en(mem_196_3_R0_en),
    .W0_addr(mem_196_3_W0_addr),
    .W0_clk(mem_196_3_W0_clk),
    .W0_data(mem_196_3_W0_data),
    .W0_en(mem_196_3_W0_en),
    .W0_mask(mem_196_3_W0_mask)
  );
  split_mem_0_ext mem_196_4 (
    .R0_addr(mem_196_4_R0_addr),
    .R0_clk(mem_196_4_R0_clk),
    .R0_data(mem_196_4_R0_data),
    .R0_en(mem_196_4_R0_en),
    .W0_addr(mem_196_4_W0_addr),
    .W0_clk(mem_196_4_W0_clk),
    .W0_data(mem_196_4_W0_data),
    .W0_en(mem_196_4_W0_en),
    .W0_mask(mem_196_4_W0_mask)
  );
  split_mem_0_ext mem_196_5 (
    .R0_addr(mem_196_5_R0_addr),
    .R0_clk(mem_196_5_R0_clk),
    .R0_data(mem_196_5_R0_data),
    .R0_en(mem_196_5_R0_en),
    .W0_addr(mem_196_5_W0_addr),
    .W0_clk(mem_196_5_W0_clk),
    .W0_data(mem_196_5_W0_data),
    .W0_en(mem_196_5_W0_en),
    .W0_mask(mem_196_5_W0_mask)
  );
  split_mem_0_ext mem_196_6 (
    .R0_addr(mem_196_6_R0_addr),
    .R0_clk(mem_196_6_R0_clk),
    .R0_data(mem_196_6_R0_data),
    .R0_en(mem_196_6_R0_en),
    .W0_addr(mem_196_6_W0_addr),
    .W0_clk(mem_196_6_W0_clk),
    .W0_data(mem_196_6_W0_data),
    .W0_en(mem_196_6_W0_en),
    .W0_mask(mem_196_6_W0_mask)
  );
  split_mem_0_ext mem_196_7 (
    .R0_addr(mem_196_7_R0_addr),
    .R0_clk(mem_196_7_R0_clk),
    .R0_data(mem_196_7_R0_data),
    .R0_en(mem_196_7_R0_en),
    .W0_addr(mem_196_7_W0_addr),
    .W0_clk(mem_196_7_W0_clk),
    .W0_data(mem_196_7_W0_data),
    .W0_en(mem_196_7_W0_en),
    .W0_mask(mem_196_7_W0_mask)
  );
  split_mem_0_ext mem_197_0 (
    .R0_addr(mem_197_0_R0_addr),
    .R0_clk(mem_197_0_R0_clk),
    .R0_data(mem_197_0_R0_data),
    .R0_en(mem_197_0_R0_en),
    .W0_addr(mem_197_0_W0_addr),
    .W0_clk(mem_197_0_W0_clk),
    .W0_data(mem_197_0_W0_data),
    .W0_en(mem_197_0_W0_en),
    .W0_mask(mem_197_0_W0_mask)
  );
  split_mem_0_ext mem_197_1 (
    .R0_addr(mem_197_1_R0_addr),
    .R0_clk(mem_197_1_R0_clk),
    .R0_data(mem_197_1_R0_data),
    .R0_en(mem_197_1_R0_en),
    .W0_addr(mem_197_1_W0_addr),
    .W0_clk(mem_197_1_W0_clk),
    .W0_data(mem_197_1_W0_data),
    .W0_en(mem_197_1_W0_en),
    .W0_mask(mem_197_1_W0_mask)
  );
  split_mem_0_ext mem_197_2 (
    .R0_addr(mem_197_2_R0_addr),
    .R0_clk(mem_197_2_R0_clk),
    .R0_data(mem_197_2_R0_data),
    .R0_en(mem_197_2_R0_en),
    .W0_addr(mem_197_2_W0_addr),
    .W0_clk(mem_197_2_W0_clk),
    .W0_data(mem_197_2_W0_data),
    .W0_en(mem_197_2_W0_en),
    .W0_mask(mem_197_2_W0_mask)
  );
  split_mem_0_ext mem_197_3 (
    .R0_addr(mem_197_3_R0_addr),
    .R0_clk(mem_197_3_R0_clk),
    .R0_data(mem_197_3_R0_data),
    .R0_en(mem_197_3_R0_en),
    .W0_addr(mem_197_3_W0_addr),
    .W0_clk(mem_197_3_W0_clk),
    .W0_data(mem_197_3_W0_data),
    .W0_en(mem_197_3_W0_en),
    .W0_mask(mem_197_3_W0_mask)
  );
  split_mem_0_ext mem_197_4 (
    .R0_addr(mem_197_4_R0_addr),
    .R0_clk(mem_197_4_R0_clk),
    .R0_data(mem_197_4_R0_data),
    .R0_en(mem_197_4_R0_en),
    .W0_addr(mem_197_4_W0_addr),
    .W0_clk(mem_197_4_W0_clk),
    .W0_data(mem_197_4_W0_data),
    .W0_en(mem_197_4_W0_en),
    .W0_mask(mem_197_4_W0_mask)
  );
  split_mem_0_ext mem_197_5 (
    .R0_addr(mem_197_5_R0_addr),
    .R0_clk(mem_197_5_R0_clk),
    .R0_data(mem_197_5_R0_data),
    .R0_en(mem_197_5_R0_en),
    .W0_addr(mem_197_5_W0_addr),
    .W0_clk(mem_197_5_W0_clk),
    .W0_data(mem_197_5_W0_data),
    .W0_en(mem_197_5_W0_en),
    .W0_mask(mem_197_5_W0_mask)
  );
  split_mem_0_ext mem_197_6 (
    .R0_addr(mem_197_6_R0_addr),
    .R0_clk(mem_197_6_R0_clk),
    .R0_data(mem_197_6_R0_data),
    .R0_en(mem_197_6_R0_en),
    .W0_addr(mem_197_6_W0_addr),
    .W0_clk(mem_197_6_W0_clk),
    .W0_data(mem_197_6_W0_data),
    .W0_en(mem_197_6_W0_en),
    .W0_mask(mem_197_6_W0_mask)
  );
  split_mem_0_ext mem_197_7 (
    .R0_addr(mem_197_7_R0_addr),
    .R0_clk(mem_197_7_R0_clk),
    .R0_data(mem_197_7_R0_data),
    .R0_en(mem_197_7_R0_en),
    .W0_addr(mem_197_7_W0_addr),
    .W0_clk(mem_197_7_W0_clk),
    .W0_data(mem_197_7_W0_data),
    .W0_en(mem_197_7_W0_en),
    .W0_mask(mem_197_7_W0_mask)
  );
  split_mem_0_ext mem_198_0 (
    .R0_addr(mem_198_0_R0_addr),
    .R0_clk(mem_198_0_R0_clk),
    .R0_data(mem_198_0_R0_data),
    .R0_en(mem_198_0_R0_en),
    .W0_addr(mem_198_0_W0_addr),
    .W0_clk(mem_198_0_W0_clk),
    .W0_data(mem_198_0_W0_data),
    .W0_en(mem_198_0_W0_en),
    .W0_mask(mem_198_0_W0_mask)
  );
  split_mem_0_ext mem_198_1 (
    .R0_addr(mem_198_1_R0_addr),
    .R0_clk(mem_198_1_R0_clk),
    .R0_data(mem_198_1_R0_data),
    .R0_en(mem_198_1_R0_en),
    .W0_addr(mem_198_1_W0_addr),
    .W0_clk(mem_198_1_W0_clk),
    .W0_data(mem_198_1_W0_data),
    .W0_en(mem_198_1_W0_en),
    .W0_mask(mem_198_1_W0_mask)
  );
  split_mem_0_ext mem_198_2 (
    .R0_addr(mem_198_2_R0_addr),
    .R0_clk(mem_198_2_R0_clk),
    .R0_data(mem_198_2_R0_data),
    .R0_en(mem_198_2_R0_en),
    .W0_addr(mem_198_2_W0_addr),
    .W0_clk(mem_198_2_W0_clk),
    .W0_data(mem_198_2_W0_data),
    .W0_en(mem_198_2_W0_en),
    .W0_mask(mem_198_2_W0_mask)
  );
  split_mem_0_ext mem_198_3 (
    .R0_addr(mem_198_3_R0_addr),
    .R0_clk(mem_198_3_R0_clk),
    .R0_data(mem_198_3_R0_data),
    .R0_en(mem_198_3_R0_en),
    .W0_addr(mem_198_3_W0_addr),
    .W0_clk(mem_198_3_W0_clk),
    .W0_data(mem_198_3_W0_data),
    .W0_en(mem_198_3_W0_en),
    .W0_mask(mem_198_3_W0_mask)
  );
  split_mem_0_ext mem_198_4 (
    .R0_addr(mem_198_4_R0_addr),
    .R0_clk(mem_198_4_R0_clk),
    .R0_data(mem_198_4_R0_data),
    .R0_en(mem_198_4_R0_en),
    .W0_addr(mem_198_4_W0_addr),
    .W0_clk(mem_198_4_W0_clk),
    .W0_data(mem_198_4_W0_data),
    .W0_en(mem_198_4_W0_en),
    .W0_mask(mem_198_4_W0_mask)
  );
  split_mem_0_ext mem_198_5 (
    .R0_addr(mem_198_5_R0_addr),
    .R0_clk(mem_198_5_R0_clk),
    .R0_data(mem_198_5_R0_data),
    .R0_en(mem_198_5_R0_en),
    .W0_addr(mem_198_5_W0_addr),
    .W0_clk(mem_198_5_W0_clk),
    .W0_data(mem_198_5_W0_data),
    .W0_en(mem_198_5_W0_en),
    .W0_mask(mem_198_5_W0_mask)
  );
  split_mem_0_ext mem_198_6 (
    .R0_addr(mem_198_6_R0_addr),
    .R0_clk(mem_198_6_R0_clk),
    .R0_data(mem_198_6_R0_data),
    .R0_en(mem_198_6_R0_en),
    .W0_addr(mem_198_6_W0_addr),
    .W0_clk(mem_198_6_W0_clk),
    .W0_data(mem_198_6_W0_data),
    .W0_en(mem_198_6_W0_en),
    .W0_mask(mem_198_6_W0_mask)
  );
  split_mem_0_ext mem_198_7 (
    .R0_addr(mem_198_7_R0_addr),
    .R0_clk(mem_198_7_R0_clk),
    .R0_data(mem_198_7_R0_data),
    .R0_en(mem_198_7_R0_en),
    .W0_addr(mem_198_7_W0_addr),
    .W0_clk(mem_198_7_W0_clk),
    .W0_data(mem_198_7_W0_data),
    .W0_en(mem_198_7_W0_en),
    .W0_mask(mem_198_7_W0_mask)
  );
  split_mem_0_ext mem_199_0 (
    .R0_addr(mem_199_0_R0_addr),
    .R0_clk(mem_199_0_R0_clk),
    .R0_data(mem_199_0_R0_data),
    .R0_en(mem_199_0_R0_en),
    .W0_addr(mem_199_0_W0_addr),
    .W0_clk(mem_199_0_W0_clk),
    .W0_data(mem_199_0_W0_data),
    .W0_en(mem_199_0_W0_en),
    .W0_mask(mem_199_0_W0_mask)
  );
  split_mem_0_ext mem_199_1 (
    .R0_addr(mem_199_1_R0_addr),
    .R0_clk(mem_199_1_R0_clk),
    .R0_data(mem_199_1_R0_data),
    .R0_en(mem_199_1_R0_en),
    .W0_addr(mem_199_1_W0_addr),
    .W0_clk(mem_199_1_W0_clk),
    .W0_data(mem_199_1_W0_data),
    .W0_en(mem_199_1_W0_en),
    .W0_mask(mem_199_1_W0_mask)
  );
  split_mem_0_ext mem_199_2 (
    .R0_addr(mem_199_2_R0_addr),
    .R0_clk(mem_199_2_R0_clk),
    .R0_data(mem_199_2_R0_data),
    .R0_en(mem_199_2_R0_en),
    .W0_addr(mem_199_2_W0_addr),
    .W0_clk(mem_199_2_W0_clk),
    .W0_data(mem_199_2_W0_data),
    .W0_en(mem_199_2_W0_en),
    .W0_mask(mem_199_2_W0_mask)
  );
  split_mem_0_ext mem_199_3 (
    .R0_addr(mem_199_3_R0_addr),
    .R0_clk(mem_199_3_R0_clk),
    .R0_data(mem_199_3_R0_data),
    .R0_en(mem_199_3_R0_en),
    .W0_addr(mem_199_3_W0_addr),
    .W0_clk(mem_199_3_W0_clk),
    .W0_data(mem_199_3_W0_data),
    .W0_en(mem_199_3_W0_en),
    .W0_mask(mem_199_3_W0_mask)
  );
  split_mem_0_ext mem_199_4 (
    .R0_addr(mem_199_4_R0_addr),
    .R0_clk(mem_199_4_R0_clk),
    .R0_data(mem_199_4_R0_data),
    .R0_en(mem_199_4_R0_en),
    .W0_addr(mem_199_4_W0_addr),
    .W0_clk(mem_199_4_W0_clk),
    .W0_data(mem_199_4_W0_data),
    .W0_en(mem_199_4_W0_en),
    .W0_mask(mem_199_4_W0_mask)
  );
  split_mem_0_ext mem_199_5 (
    .R0_addr(mem_199_5_R0_addr),
    .R0_clk(mem_199_5_R0_clk),
    .R0_data(mem_199_5_R0_data),
    .R0_en(mem_199_5_R0_en),
    .W0_addr(mem_199_5_W0_addr),
    .W0_clk(mem_199_5_W0_clk),
    .W0_data(mem_199_5_W0_data),
    .W0_en(mem_199_5_W0_en),
    .W0_mask(mem_199_5_W0_mask)
  );
  split_mem_0_ext mem_199_6 (
    .R0_addr(mem_199_6_R0_addr),
    .R0_clk(mem_199_6_R0_clk),
    .R0_data(mem_199_6_R0_data),
    .R0_en(mem_199_6_R0_en),
    .W0_addr(mem_199_6_W0_addr),
    .W0_clk(mem_199_6_W0_clk),
    .W0_data(mem_199_6_W0_data),
    .W0_en(mem_199_6_W0_en),
    .W0_mask(mem_199_6_W0_mask)
  );
  split_mem_0_ext mem_199_7 (
    .R0_addr(mem_199_7_R0_addr),
    .R0_clk(mem_199_7_R0_clk),
    .R0_data(mem_199_7_R0_data),
    .R0_en(mem_199_7_R0_en),
    .W0_addr(mem_199_7_W0_addr),
    .W0_clk(mem_199_7_W0_clk),
    .W0_data(mem_199_7_W0_data),
    .W0_en(mem_199_7_W0_en),
    .W0_mask(mem_199_7_W0_mask)
  );
  split_mem_0_ext mem_200_0 (
    .R0_addr(mem_200_0_R0_addr),
    .R0_clk(mem_200_0_R0_clk),
    .R0_data(mem_200_0_R0_data),
    .R0_en(mem_200_0_R0_en),
    .W0_addr(mem_200_0_W0_addr),
    .W0_clk(mem_200_0_W0_clk),
    .W0_data(mem_200_0_W0_data),
    .W0_en(mem_200_0_W0_en),
    .W0_mask(mem_200_0_W0_mask)
  );
  split_mem_0_ext mem_200_1 (
    .R0_addr(mem_200_1_R0_addr),
    .R0_clk(mem_200_1_R0_clk),
    .R0_data(mem_200_1_R0_data),
    .R0_en(mem_200_1_R0_en),
    .W0_addr(mem_200_1_W0_addr),
    .W0_clk(mem_200_1_W0_clk),
    .W0_data(mem_200_1_W0_data),
    .W0_en(mem_200_1_W0_en),
    .W0_mask(mem_200_1_W0_mask)
  );
  split_mem_0_ext mem_200_2 (
    .R0_addr(mem_200_2_R0_addr),
    .R0_clk(mem_200_2_R0_clk),
    .R0_data(mem_200_2_R0_data),
    .R0_en(mem_200_2_R0_en),
    .W0_addr(mem_200_2_W0_addr),
    .W0_clk(mem_200_2_W0_clk),
    .W0_data(mem_200_2_W0_data),
    .W0_en(mem_200_2_W0_en),
    .W0_mask(mem_200_2_W0_mask)
  );
  split_mem_0_ext mem_200_3 (
    .R0_addr(mem_200_3_R0_addr),
    .R0_clk(mem_200_3_R0_clk),
    .R0_data(mem_200_3_R0_data),
    .R0_en(mem_200_3_R0_en),
    .W0_addr(mem_200_3_W0_addr),
    .W0_clk(mem_200_3_W0_clk),
    .W0_data(mem_200_3_W0_data),
    .W0_en(mem_200_3_W0_en),
    .W0_mask(mem_200_3_W0_mask)
  );
  split_mem_0_ext mem_200_4 (
    .R0_addr(mem_200_4_R0_addr),
    .R0_clk(mem_200_4_R0_clk),
    .R0_data(mem_200_4_R0_data),
    .R0_en(mem_200_4_R0_en),
    .W0_addr(mem_200_4_W0_addr),
    .W0_clk(mem_200_4_W0_clk),
    .W0_data(mem_200_4_W0_data),
    .W0_en(mem_200_4_W0_en),
    .W0_mask(mem_200_4_W0_mask)
  );
  split_mem_0_ext mem_200_5 (
    .R0_addr(mem_200_5_R0_addr),
    .R0_clk(mem_200_5_R0_clk),
    .R0_data(mem_200_5_R0_data),
    .R0_en(mem_200_5_R0_en),
    .W0_addr(mem_200_5_W0_addr),
    .W0_clk(mem_200_5_W0_clk),
    .W0_data(mem_200_5_W0_data),
    .W0_en(mem_200_5_W0_en),
    .W0_mask(mem_200_5_W0_mask)
  );
  split_mem_0_ext mem_200_6 (
    .R0_addr(mem_200_6_R0_addr),
    .R0_clk(mem_200_6_R0_clk),
    .R0_data(mem_200_6_R0_data),
    .R0_en(mem_200_6_R0_en),
    .W0_addr(mem_200_6_W0_addr),
    .W0_clk(mem_200_6_W0_clk),
    .W0_data(mem_200_6_W0_data),
    .W0_en(mem_200_6_W0_en),
    .W0_mask(mem_200_6_W0_mask)
  );
  split_mem_0_ext mem_200_7 (
    .R0_addr(mem_200_7_R0_addr),
    .R0_clk(mem_200_7_R0_clk),
    .R0_data(mem_200_7_R0_data),
    .R0_en(mem_200_7_R0_en),
    .W0_addr(mem_200_7_W0_addr),
    .W0_clk(mem_200_7_W0_clk),
    .W0_data(mem_200_7_W0_data),
    .W0_en(mem_200_7_W0_en),
    .W0_mask(mem_200_7_W0_mask)
  );
  split_mem_0_ext mem_201_0 (
    .R0_addr(mem_201_0_R0_addr),
    .R0_clk(mem_201_0_R0_clk),
    .R0_data(mem_201_0_R0_data),
    .R0_en(mem_201_0_R0_en),
    .W0_addr(mem_201_0_W0_addr),
    .W0_clk(mem_201_0_W0_clk),
    .W0_data(mem_201_0_W0_data),
    .W0_en(mem_201_0_W0_en),
    .W0_mask(mem_201_0_W0_mask)
  );
  split_mem_0_ext mem_201_1 (
    .R0_addr(mem_201_1_R0_addr),
    .R0_clk(mem_201_1_R0_clk),
    .R0_data(mem_201_1_R0_data),
    .R0_en(mem_201_1_R0_en),
    .W0_addr(mem_201_1_W0_addr),
    .W0_clk(mem_201_1_W0_clk),
    .W0_data(mem_201_1_W0_data),
    .W0_en(mem_201_1_W0_en),
    .W0_mask(mem_201_1_W0_mask)
  );
  split_mem_0_ext mem_201_2 (
    .R0_addr(mem_201_2_R0_addr),
    .R0_clk(mem_201_2_R0_clk),
    .R0_data(mem_201_2_R0_data),
    .R0_en(mem_201_2_R0_en),
    .W0_addr(mem_201_2_W0_addr),
    .W0_clk(mem_201_2_W0_clk),
    .W0_data(mem_201_2_W0_data),
    .W0_en(mem_201_2_W0_en),
    .W0_mask(mem_201_2_W0_mask)
  );
  split_mem_0_ext mem_201_3 (
    .R0_addr(mem_201_3_R0_addr),
    .R0_clk(mem_201_3_R0_clk),
    .R0_data(mem_201_3_R0_data),
    .R0_en(mem_201_3_R0_en),
    .W0_addr(mem_201_3_W0_addr),
    .W0_clk(mem_201_3_W0_clk),
    .W0_data(mem_201_3_W0_data),
    .W0_en(mem_201_3_W0_en),
    .W0_mask(mem_201_3_W0_mask)
  );
  split_mem_0_ext mem_201_4 (
    .R0_addr(mem_201_4_R0_addr),
    .R0_clk(mem_201_4_R0_clk),
    .R0_data(mem_201_4_R0_data),
    .R0_en(mem_201_4_R0_en),
    .W0_addr(mem_201_4_W0_addr),
    .W0_clk(mem_201_4_W0_clk),
    .W0_data(mem_201_4_W0_data),
    .W0_en(mem_201_4_W0_en),
    .W0_mask(mem_201_4_W0_mask)
  );
  split_mem_0_ext mem_201_5 (
    .R0_addr(mem_201_5_R0_addr),
    .R0_clk(mem_201_5_R0_clk),
    .R0_data(mem_201_5_R0_data),
    .R0_en(mem_201_5_R0_en),
    .W0_addr(mem_201_5_W0_addr),
    .W0_clk(mem_201_5_W0_clk),
    .W0_data(mem_201_5_W0_data),
    .W0_en(mem_201_5_W0_en),
    .W0_mask(mem_201_5_W0_mask)
  );
  split_mem_0_ext mem_201_6 (
    .R0_addr(mem_201_6_R0_addr),
    .R0_clk(mem_201_6_R0_clk),
    .R0_data(mem_201_6_R0_data),
    .R0_en(mem_201_6_R0_en),
    .W0_addr(mem_201_6_W0_addr),
    .W0_clk(mem_201_6_W0_clk),
    .W0_data(mem_201_6_W0_data),
    .W0_en(mem_201_6_W0_en),
    .W0_mask(mem_201_6_W0_mask)
  );
  split_mem_0_ext mem_201_7 (
    .R0_addr(mem_201_7_R0_addr),
    .R0_clk(mem_201_7_R0_clk),
    .R0_data(mem_201_7_R0_data),
    .R0_en(mem_201_7_R0_en),
    .W0_addr(mem_201_7_W0_addr),
    .W0_clk(mem_201_7_W0_clk),
    .W0_data(mem_201_7_W0_data),
    .W0_en(mem_201_7_W0_en),
    .W0_mask(mem_201_7_W0_mask)
  );
  split_mem_0_ext mem_202_0 (
    .R0_addr(mem_202_0_R0_addr),
    .R0_clk(mem_202_0_R0_clk),
    .R0_data(mem_202_0_R0_data),
    .R0_en(mem_202_0_R0_en),
    .W0_addr(mem_202_0_W0_addr),
    .W0_clk(mem_202_0_W0_clk),
    .W0_data(mem_202_0_W0_data),
    .W0_en(mem_202_0_W0_en),
    .W0_mask(mem_202_0_W0_mask)
  );
  split_mem_0_ext mem_202_1 (
    .R0_addr(mem_202_1_R0_addr),
    .R0_clk(mem_202_1_R0_clk),
    .R0_data(mem_202_1_R0_data),
    .R0_en(mem_202_1_R0_en),
    .W0_addr(mem_202_1_W0_addr),
    .W0_clk(mem_202_1_W0_clk),
    .W0_data(mem_202_1_W0_data),
    .W0_en(mem_202_1_W0_en),
    .W0_mask(mem_202_1_W0_mask)
  );
  split_mem_0_ext mem_202_2 (
    .R0_addr(mem_202_2_R0_addr),
    .R0_clk(mem_202_2_R0_clk),
    .R0_data(mem_202_2_R0_data),
    .R0_en(mem_202_2_R0_en),
    .W0_addr(mem_202_2_W0_addr),
    .W0_clk(mem_202_2_W0_clk),
    .W0_data(mem_202_2_W0_data),
    .W0_en(mem_202_2_W0_en),
    .W0_mask(mem_202_2_W0_mask)
  );
  split_mem_0_ext mem_202_3 (
    .R0_addr(mem_202_3_R0_addr),
    .R0_clk(mem_202_3_R0_clk),
    .R0_data(mem_202_3_R0_data),
    .R0_en(mem_202_3_R0_en),
    .W0_addr(mem_202_3_W0_addr),
    .W0_clk(mem_202_3_W0_clk),
    .W0_data(mem_202_3_W0_data),
    .W0_en(mem_202_3_W0_en),
    .W0_mask(mem_202_3_W0_mask)
  );
  split_mem_0_ext mem_202_4 (
    .R0_addr(mem_202_4_R0_addr),
    .R0_clk(mem_202_4_R0_clk),
    .R0_data(mem_202_4_R0_data),
    .R0_en(mem_202_4_R0_en),
    .W0_addr(mem_202_4_W0_addr),
    .W0_clk(mem_202_4_W0_clk),
    .W0_data(mem_202_4_W0_data),
    .W0_en(mem_202_4_W0_en),
    .W0_mask(mem_202_4_W0_mask)
  );
  split_mem_0_ext mem_202_5 (
    .R0_addr(mem_202_5_R0_addr),
    .R0_clk(mem_202_5_R0_clk),
    .R0_data(mem_202_5_R0_data),
    .R0_en(mem_202_5_R0_en),
    .W0_addr(mem_202_5_W0_addr),
    .W0_clk(mem_202_5_W0_clk),
    .W0_data(mem_202_5_W0_data),
    .W0_en(mem_202_5_W0_en),
    .W0_mask(mem_202_5_W0_mask)
  );
  split_mem_0_ext mem_202_6 (
    .R0_addr(mem_202_6_R0_addr),
    .R0_clk(mem_202_6_R0_clk),
    .R0_data(mem_202_6_R0_data),
    .R0_en(mem_202_6_R0_en),
    .W0_addr(mem_202_6_W0_addr),
    .W0_clk(mem_202_6_W0_clk),
    .W0_data(mem_202_6_W0_data),
    .W0_en(mem_202_6_W0_en),
    .W0_mask(mem_202_6_W0_mask)
  );
  split_mem_0_ext mem_202_7 (
    .R0_addr(mem_202_7_R0_addr),
    .R0_clk(mem_202_7_R0_clk),
    .R0_data(mem_202_7_R0_data),
    .R0_en(mem_202_7_R0_en),
    .W0_addr(mem_202_7_W0_addr),
    .W0_clk(mem_202_7_W0_clk),
    .W0_data(mem_202_7_W0_data),
    .W0_en(mem_202_7_W0_en),
    .W0_mask(mem_202_7_W0_mask)
  );
  split_mem_0_ext mem_203_0 (
    .R0_addr(mem_203_0_R0_addr),
    .R0_clk(mem_203_0_R0_clk),
    .R0_data(mem_203_0_R0_data),
    .R0_en(mem_203_0_R0_en),
    .W0_addr(mem_203_0_W0_addr),
    .W0_clk(mem_203_0_W0_clk),
    .W0_data(mem_203_0_W0_data),
    .W0_en(mem_203_0_W0_en),
    .W0_mask(mem_203_0_W0_mask)
  );
  split_mem_0_ext mem_203_1 (
    .R0_addr(mem_203_1_R0_addr),
    .R0_clk(mem_203_1_R0_clk),
    .R0_data(mem_203_1_R0_data),
    .R0_en(mem_203_1_R0_en),
    .W0_addr(mem_203_1_W0_addr),
    .W0_clk(mem_203_1_W0_clk),
    .W0_data(mem_203_1_W0_data),
    .W0_en(mem_203_1_W0_en),
    .W0_mask(mem_203_1_W0_mask)
  );
  split_mem_0_ext mem_203_2 (
    .R0_addr(mem_203_2_R0_addr),
    .R0_clk(mem_203_2_R0_clk),
    .R0_data(mem_203_2_R0_data),
    .R0_en(mem_203_2_R0_en),
    .W0_addr(mem_203_2_W0_addr),
    .W0_clk(mem_203_2_W0_clk),
    .W0_data(mem_203_2_W0_data),
    .W0_en(mem_203_2_W0_en),
    .W0_mask(mem_203_2_W0_mask)
  );
  split_mem_0_ext mem_203_3 (
    .R0_addr(mem_203_3_R0_addr),
    .R0_clk(mem_203_3_R0_clk),
    .R0_data(mem_203_3_R0_data),
    .R0_en(mem_203_3_R0_en),
    .W0_addr(mem_203_3_W0_addr),
    .W0_clk(mem_203_3_W0_clk),
    .W0_data(mem_203_3_W0_data),
    .W0_en(mem_203_3_W0_en),
    .W0_mask(mem_203_3_W0_mask)
  );
  split_mem_0_ext mem_203_4 (
    .R0_addr(mem_203_4_R0_addr),
    .R0_clk(mem_203_4_R0_clk),
    .R0_data(mem_203_4_R0_data),
    .R0_en(mem_203_4_R0_en),
    .W0_addr(mem_203_4_W0_addr),
    .W0_clk(mem_203_4_W0_clk),
    .W0_data(mem_203_4_W0_data),
    .W0_en(mem_203_4_W0_en),
    .W0_mask(mem_203_4_W0_mask)
  );
  split_mem_0_ext mem_203_5 (
    .R0_addr(mem_203_5_R0_addr),
    .R0_clk(mem_203_5_R0_clk),
    .R0_data(mem_203_5_R0_data),
    .R0_en(mem_203_5_R0_en),
    .W0_addr(mem_203_5_W0_addr),
    .W0_clk(mem_203_5_W0_clk),
    .W0_data(mem_203_5_W0_data),
    .W0_en(mem_203_5_W0_en),
    .W0_mask(mem_203_5_W0_mask)
  );
  split_mem_0_ext mem_203_6 (
    .R0_addr(mem_203_6_R0_addr),
    .R0_clk(mem_203_6_R0_clk),
    .R0_data(mem_203_6_R0_data),
    .R0_en(mem_203_6_R0_en),
    .W0_addr(mem_203_6_W0_addr),
    .W0_clk(mem_203_6_W0_clk),
    .W0_data(mem_203_6_W0_data),
    .W0_en(mem_203_6_W0_en),
    .W0_mask(mem_203_6_W0_mask)
  );
  split_mem_0_ext mem_203_7 (
    .R0_addr(mem_203_7_R0_addr),
    .R0_clk(mem_203_7_R0_clk),
    .R0_data(mem_203_7_R0_data),
    .R0_en(mem_203_7_R0_en),
    .W0_addr(mem_203_7_W0_addr),
    .W0_clk(mem_203_7_W0_clk),
    .W0_data(mem_203_7_W0_data),
    .W0_en(mem_203_7_W0_en),
    .W0_mask(mem_203_7_W0_mask)
  );
  split_mem_0_ext mem_204_0 (
    .R0_addr(mem_204_0_R0_addr),
    .R0_clk(mem_204_0_R0_clk),
    .R0_data(mem_204_0_R0_data),
    .R0_en(mem_204_0_R0_en),
    .W0_addr(mem_204_0_W0_addr),
    .W0_clk(mem_204_0_W0_clk),
    .W0_data(mem_204_0_W0_data),
    .W0_en(mem_204_0_W0_en),
    .W0_mask(mem_204_0_W0_mask)
  );
  split_mem_0_ext mem_204_1 (
    .R0_addr(mem_204_1_R0_addr),
    .R0_clk(mem_204_1_R0_clk),
    .R0_data(mem_204_1_R0_data),
    .R0_en(mem_204_1_R0_en),
    .W0_addr(mem_204_1_W0_addr),
    .W0_clk(mem_204_1_W0_clk),
    .W0_data(mem_204_1_W0_data),
    .W0_en(mem_204_1_W0_en),
    .W0_mask(mem_204_1_W0_mask)
  );
  split_mem_0_ext mem_204_2 (
    .R0_addr(mem_204_2_R0_addr),
    .R0_clk(mem_204_2_R0_clk),
    .R0_data(mem_204_2_R0_data),
    .R0_en(mem_204_2_R0_en),
    .W0_addr(mem_204_2_W0_addr),
    .W0_clk(mem_204_2_W0_clk),
    .W0_data(mem_204_2_W0_data),
    .W0_en(mem_204_2_W0_en),
    .W0_mask(mem_204_2_W0_mask)
  );
  split_mem_0_ext mem_204_3 (
    .R0_addr(mem_204_3_R0_addr),
    .R0_clk(mem_204_3_R0_clk),
    .R0_data(mem_204_3_R0_data),
    .R0_en(mem_204_3_R0_en),
    .W0_addr(mem_204_3_W0_addr),
    .W0_clk(mem_204_3_W0_clk),
    .W0_data(mem_204_3_W0_data),
    .W0_en(mem_204_3_W0_en),
    .W0_mask(mem_204_3_W0_mask)
  );
  split_mem_0_ext mem_204_4 (
    .R0_addr(mem_204_4_R0_addr),
    .R0_clk(mem_204_4_R0_clk),
    .R0_data(mem_204_4_R0_data),
    .R0_en(mem_204_4_R0_en),
    .W0_addr(mem_204_4_W0_addr),
    .W0_clk(mem_204_4_W0_clk),
    .W0_data(mem_204_4_W0_data),
    .W0_en(mem_204_4_W0_en),
    .W0_mask(mem_204_4_W0_mask)
  );
  split_mem_0_ext mem_204_5 (
    .R0_addr(mem_204_5_R0_addr),
    .R0_clk(mem_204_5_R0_clk),
    .R0_data(mem_204_5_R0_data),
    .R0_en(mem_204_5_R0_en),
    .W0_addr(mem_204_5_W0_addr),
    .W0_clk(mem_204_5_W0_clk),
    .W0_data(mem_204_5_W0_data),
    .W0_en(mem_204_5_W0_en),
    .W0_mask(mem_204_5_W0_mask)
  );
  split_mem_0_ext mem_204_6 (
    .R0_addr(mem_204_6_R0_addr),
    .R0_clk(mem_204_6_R0_clk),
    .R0_data(mem_204_6_R0_data),
    .R0_en(mem_204_6_R0_en),
    .W0_addr(mem_204_6_W0_addr),
    .W0_clk(mem_204_6_W0_clk),
    .W0_data(mem_204_6_W0_data),
    .W0_en(mem_204_6_W0_en),
    .W0_mask(mem_204_6_W0_mask)
  );
  split_mem_0_ext mem_204_7 (
    .R0_addr(mem_204_7_R0_addr),
    .R0_clk(mem_204_7_R0_clk),
    .R0_data(mem_204_7_R0_data),
    .R0_en(mem_204_7_R0_en),
    .W0_addr(mem_204_7_W0_addr),
    .W0_clk(mem_204_7_W0_clk),
    .W0_data(mem_204_7_W0_data),
    .W0_en(mem_204_7_W0_en),
    .W0_mask(mem_204_7_W0_mask)
  );
  split_mem_0_ext mem_205_0 (
    .R0_addr(mem_205_0_R0_addr),
    .R0_clk(mem_205_0_R0_clk),
    .R0_data(mem_205_0_R0_data),
    .R0_en(mem_205_0_R0_en),
    .W0_addr(mem_205_0_W0_addr),
    .W0_clk(mem_205_0_W0_clk),
    .W0_data(mem_205_0_W0_data),
    .W0_en(mem_205_0_W0_en),
    .W0_mask(mem_205_0_W0_mask)
  );
  split_mem_0_ext mem_205_1 (
    .R0_addr(mem_205_1_R0_addr),
    .R0_clk(mem_205_1_R0_clk),
    .R0_data(mem_205_1_R0_data),
    .R0_en(mem_205_1_R0_en),
    .W0_addr(mem_205_1_W0_addr),
    .W0_clk(mem_205_1_W0_clk),
    .W0_data(mem_205_1_W0_data),
    .W0_en(mem_205_1_W0_en),
    .W0_mask(mem_205_1_W0_mask)
  );
  split_mem_0_ext mem_205_2 (
    .R0_addr(mem_205_2_R0_addr),
    .R0_clk(mem_205_2_R0_clk),
    .R0_data(mem_205_2_R0_data),
    .R0_en(mem_205_2_R0_en),
    .W0_addr(mem_205_2_W0_addr),
    .W0_clk(mem_205_2_W0_clk),
    .W0_data(mem_205_2_W0_data),
    .W0_en(mem_205_2_W0_en),
    .W0_mask(mem_205_2_W0_mask)
  );
  split_mem_0_ext mem_205_3 (
    .R0_addr(mem_205_3_R0_addr),
    .R0_clk(mem_205_3_R0_clk),
    .R0_data(mem_205_3_R0_data),
    .R0_en(mem_205_3_R0_en),
    .W0_addr(mem_205_3_W0_addr),
    .W0_clk(mem_205_3_W0_clk),
    .W0_data(mem_205_3_W0_data),
    .W0_en(mem_205_3_W0_en),
    .W0_mask(mem_205_3_W0_mask)
  );
  split_mem_0_ext mem_205_4 (
    .R0_addr(mem_205_4_R0_addr),
    .R0_clk(mem_205_4_R0_clk),
    .R0_data(mem_205_4_R0_data),
    .R0_en(mem_205_4_R0_en),
    .W0_addr(mem_205_4_W0_addr),
    .W0_clk(mem_205_4_W0_clk),
    .W0_data(mem_205_4_W0_data),
    .W0_en(mem_205_4_W0_en),
    .W0_mask(mem_205_4_W0_mask)
  );
  split_mem_0_ext mem_205_5 (
    .R0_addr(mem_205_5_R0_addr),
    .R0_clk(mem_205_5_R0_clk),
    .R0_data(mem_205_5_R0_data),
    .R0_en(mem_205_5_R0_en),
    .W0_addr(mem_205_5_W0_addr),
    .W0_clk(mem_205_5_W0_clk),
    .W0_data(mem_205_5_W0_data),
    .W0_en(mem_205_5_W0_en),
    .W0_mask(mem_205_5_W0_mask)
  );
  split_mem_0_ext mem_205_6 (
    .R0_addr(mem_205_6_R0_addr),
    .R0_clk(mem_205_6_R0_clk),
    .R0_data(mem_205_6_R0_data),
    .R0_en(mem_205_6_R0_en),
    .W0_addr(mem_205_6_W0_addr),
    .W0_clk(mem_205_6_W0_clk),
    .W0_data(mem_205_6_W0_data),
    .W0_en(mem_205_6_W0_en),
    .W0_mask(mem_205_6_W0_mask)
  );
  split_mem_0_ext mem_205_7 (
    .R0_addr(mem_205_7_R0_addr),
    .R0_clk(mem_205_7_R0_clk),
    .R0_data(mem_205_7_R0_data),
    .R0_en(mem_205_7_R0_en),
    .W0_addr(mem_205_7_W0_addr),
    .W0_clk(mem_205_7_W0_clk),
    .W0_data(mem_205_7_W0_data),
    .W0_en(mem_205_7_W0_en),
    .W0_mask(mem_205_7_W0_mask)
  );
  split_mem_0_ext mem_206_0 (
    .R0_addr(mem_206_0_R0_addr),
    .R0_clk(mem_206_0_R0_clk),
    .R0_data(mem_206_0_R0_data),
    .R0_en(mem_206_0_R0_en),
    .W0_addr(mem_206_0_W0_addr),
    .W0_clk(mem_206_0_W0_clk),
    .W0_data(mem_206_0_W0_data),
    .W0_en(mem_206_0_W0_en),
    .W0_mask(mem_206_0_W0_mask)
  );
  split_mem_0_ext mem_206_1 (
    .R0_addr(mem_206_1_R0_addr),
    .R0_clk(mem_206_1_R0_clk),
    .R0_data(mem_206_1_R0_data),
    .R0_en(mem_206_1_R0_en),
    .W0_addr(mem_206_1_W0_addr),
    .W0_clk(mem_206_1_W0_clk),
    .W0_data(mem_206_1_W0_data),
    .W0_en(mem_206_1_W0_en),
    .W0_mask(mem_206_1_W0_mask)
  );
  split_mem_0_ext mem_206_2 (
    .R0_addr(mem_206_2_R0_addr),
    .R0_clk(mem_206_2_R0_clk),
    .R0_data(mem_206_2_R0_data),
    .R0_en(mem_206_2_R0_en),
    .W0_addr(mem_206_2_W0_addr),
    .W0_clk(mem_206_2_W0_clk),
    .W0_data(mem_206_2_W0_data),
    .W0_en(mem_206_2_W0_en),
    .W0_mask(mem_206_2_W0_mask)
  );
  split_mem_0_ext mem_206_3 (
    .R0_addr(mem_206_3_R0_addr),
    .R0_clk(mem_206_3_R0_clk),
    .R0_data(mem_206_3_R0_data),
    .R0_en(mem_206_3_R0_en),
    .W0_addr(mem_206_3_W0_addr),
    .W0_clk(mem_206_3_W0_clk),
    .W0_data(mem_206_3_W0_data),
    .W0_en(mem_206_3_W0_en),
    .W0_mask(mem_206_3_W0_mask)
  );
  split_mem_0_ext mem_206_4 (
    .R0_addr(mem_206_4_R0_addr),
    .R0_clk(mem_206_4_R0_clk),
    .R0_data(mem_206_4_R0_data),
    .R0_en(mem_206_4_R0_en),
    .W0_addr(mem_206_4_W0_addr),
    .W0_clk(mem_206_4_W0_clk),
    .W0_data(mem_206_4_W0_data),
    .W0_en(mem_206_4_W0_en),
    .W0_mask(mem_206_4_W0_mask)
  );
  split_mem_0_ext mem_206_5 (
    .R0_addr(mem_206_5_R0_addr),
    .R0_clk(mem_206_5_R0_clk),
    .R0_data(mem_206_5_R0_data),
    .R0_en(mem_206_5_R0_en),
    .W0_addr(mem_206_5_W0_addr),
    .W0_clk(mem_206_5_W0_clk),
    .W0_data(mem_206_5_W0_data),
    .W0_en(mem_206_5_W0_en),
    .W0_mask(mem_206_5_W0_mask)
  );
  split_mem_0_ext mem_206_6 (
    .R0_addr(mem_206_6_R0_addr),
    .R0_clk(mem_206_6_R0_clk),
    .R0_data(mem_206_6_R0_data),
    .R0_en(mem_206_6_R0_en),
    .W0_addr(mem_206_6_W0_addr),
    .W0_clk(mem_206_6_W0_clk),
    .W0_data(mem_206_6_W0_data),
    .W0_en(mem_206_6_W0_en),
    .W0_mask(mem_206_6_W0_mask)
  );
  split_mem_0_ext mem_206_7 (
    .R0_addr(mem_206_7_R0_addr),
    .R0_clk(mem_206_7_R0_clk),
    .R0_data(mem_206_7_R0_data),
    .R0_en(mem_206_7_R0_en),
    .W0_addr(mem_206_7_W0_addr),
    .W0_clk(mem_206_7_W0_clk),
    .W0_data(mem_206_7_W0_data),
    .W0_en(mem_206_7_W0_en),
    .W0_mask(mem_206_7_W0_mask)
  );
  split_mem_0_ext mem_207_0 (
    .R0_addr(mem_207_0_R0_addr),
    .R0_clk(mem_207_0_R0_clk),
    .R0_data(mem_207_0_R0_data),
    .R0_en(mem_207_0_R0_en),
    .W0_addr(mem_207_0_W0_addr),
    .W0_clk(mem_207_0_W0_clk),
    .W0_data(mem_207_0_W0_data),
    .W0_en(mem_207_0_W0_en),
    .W0_mask(mem_207_0_W0_mask)
  );
  split_mem_0_ext mem_207_1 (
    .R0_addr(mem_207_1_R0_addr),
    .R0_clk(mem_207_1_R0_clk),
    .R0_data(mem_207_1_R0_data),
    .R0_en(mem_207_1_R0_en),
    .W0_addr(mem_207_1_W0_addr),
    .W0_clk(mem_207_1_W0_clk),
    .W0_data(mem_207_1_W0_data),
    .W0_en(mem_207_1_W0_en),
    .W0_mask(mem_207_1_W0_mask)
  );
  split_mem_0_ext mem_207_2 (
    .R0_addr(mem_207_2_R0_addr),
    .R0_clk(mem_207_2_R0_clk),
    .R0_data(mem_207_2_R0_data),
    .R0_en(mem_207_2_R0_en),
    .W0_addr(mem_207_2_W0_addr),
    .W0_clk(mem_207_2_W0_clk),
    .W0_data(mem_207_2_W0_data),
    .W0_en(mem_207_2_W0_en),
    .W0_mask(mem_207_2_W0_mask)
  );
  split_mem_0_ext mem_207_3 (
    .R0_addr(mem_207_3_R0_addr),
    .R0_clk(mem_207_3_R0_clk),
    .R0_data(mem_207_3_R0_data),
    .R0_en(mem_207_3_R0_en),
    .W0_addr(mem_207_3_W0_addr),
    .W0_clk(mem_207_3_W0_clk),
    .W0_data(mem_207_3_W0_data),
    .W0_en(mem_207_3_W0_en),
    .W0_mask(mem_207_3_W0_mask)
  );
  split_mem_0_ext mem_207_4 (
    .R0_addr(mem_207_4_R0_addr),
    .R0_clk(mem_207_4_R0_clk),
    .R0_data(mem_207_4_R0_data),
    .R0_en(mem_207_4_R0_en),
    .W0_addr(mem_207_4_W0_addr),
    .W0_clk(mem_207_4_W0_clk),
    .W0_data(mem_207_4_W0_data),
    .W0_en(mem_207_4_W0_en),
    .W0_mask(mem_207_4_W0_mask)
  );
  split_mem_0_ext mem_207_5 (
    .R0_addr(mem_207_5_R0_addr),
    .R0_clk(mem_207_5_R0_clk),
    .R0_data(mem_207_5_R0_data),
    .R0_en(mem_207_5_R0_en),
    .W0_addr(mem_207_5_W0_addr),
    .W0_clk(mem_207_5_W0_clk),
    .W0_data(mem_207_5_W0_data),
    .W0_en(mem_207_5_W0_en),
    .W0_mask(mem_207_5_W0_mask)
  );
  split_mem_0_ext mem_207_6 (
    .R0_addr(mem_207_6_R0_addr),
    .R0_clk(mem_207_6_R0_clk),
    .R0_data(mem_207_6_R0_data),
    .R0_en(mem_207_6_R0_en),
    .W0_addr(mem_207_6_W0_addr),
    .W0_clk(mem_207_6_W0_clk),
    .W0_data(mem_207_6_W0_data),
    .W0_en(mem_207_6_W0_en),
    .W0_mask(mem_207_6_W0_mask)
  );
  split_mem_0_ext mem_207_7 (
    .R0_addr(mem_207_7_R0_addr),
    .R0_clk(mem_207_7_R0_clk),
    .R0_data(mem_207_7_R0_data),
    .R0_en(mem_207_7_R0_en),
    .W0_addr(mem_207_7_W0_addr),
    .W0_clk(mem_207_7_W0_clk),
    .W0_data(mem_207_7_W0_data),
    .W0_en(mem_207_7_W0_en),
    .W0_mask(mem_207_7_W0_mask)
  );
  split_mem_0_ext mem_208_0 (
    .R0_addr(mem_208_0_R0_addr),
    .R0_clk(mem_208_0_R0_clk),
    .R0_data(mem_208_0_R0_data),
    .R0_en(mem_208_0_R0_en),
    .W0_addr(mem_208_0_W0_addr),
    .W0_clk(mem_208_0_W0_clk),
    .W0_data(mem_208_0_W0_data),
    .W0_en(mem_208_0_W0_en),
    .W0_mask(mem_208_0_W0_mask)
  );
  split_mem_0_ext mem_208_1 (
    .R0_addr(mem_208_1_R0_addr),
    .R0_clk(mem_208_1_R0_clk),
    .R0_data(mem_208_1_R0_data),
    .R0_en(mem_208_1_R0_en),
    .W0_addr(mem_208_1_W0_addr),
    .W0_clk(mem_208_1_W0_clk),
    .W0_data(mem_208_1_W0_data),
    .W0_en(mem_208_1_W0_en),
    .W0_mask(mem_208_1_W0_mask)
  );
  split_mem_0_ext mem_208_2 (
    .R0_addr(mem_208_2_R0_addr),
    .R0_clk(mem_208_2_R0_clk),
    .R0_data(mem_208_2_R0_data),
    .R0_en(mem_208_2_R0_en),
    .W0_addr(mem_208_2_W0_addr),
    .W0_clk(mem_208_2_W0_clk),
    .W0_data(mem_208_2_W0_data),
    .W0_en(mem_208_2_W0_en),
    .W0_mask(mem_208_2_W0_mask)
  );
  split_mem_0_ext mem_208_3 (
    .R0_addr(mem_208_3_R0_addr),
    .R0_clk(mem_208_3_R0_clk),
    .R0_data(mem_208_3_R0_data),
    .R0_en(mem_208_3_R0_en),
    .W0_addr(mem_208_3_W0_addr),
    .W0_clk(mem_208_3_W0_clk),
    .W0_data(mem_208_3_W0_data),
    .W0_en(mem_208_3_W0_en),
    .W0_mask(mem_208_3_W0_mask)
  );
  split_mem_0_ext mem_208_4 (
    .R0_addr(mem_208_4_R0_addr),
    .R0_clk(mem_208_4_R0_clk),
    .R0_data(mem_208_4_R0_data),
    .R0_en(mem_208_4_R0_en),
    .W0_addr(mem_208_4_W0_addr),
    .W0_clk(mem_208_4_W0_clk),
    .W0_data(mem_208_4_W0_data),
    .W0_en(mem_208_4_W0_en),
    .W0_mask(mem_208_4_W0_mask)
  );
  split_mem_0_ext mem_208_5 (
    .R0_addr(mem_208_5_R0_addr),
    .R0_clk(mem_208_5_R0_clk),
    .R0_data(mem_208_5_R0_data),
    .R0_en(mem_208_5_R0_en),
    .W0_addr(mem_208_5_W0_addr),
    .W0_clk(mem_208_5_W0_clk),
    .W0_data(mem_208_5_W0_data),
    .W0_en(mem_208_5_W0_en),
    .W0_mask(mem_208_5_W0_mask)
  );
  split_mem_0_ext mem_208_6 (
    .R0_addr(mem_208_6_R0_addr),
    .R0_clk(mem_208_6_R0_clk),
    .R0_data(mem_208_6_R0_data),
    .R0_en(mem_208_6_R0_en),
    .W0_addr(mem_208_6_W0_addr),
    .W0_clk(mem_208_6_W0_clk),
    .W0_data(mem_208_6_W0_data),
    .W0_en(mem_208_6_W0_en),
    .W0_mask(mem_208_6_W0_mask)
  );
  split_mem_0_ext mem_208_7 (
    .R0_addr(mem_208_7_R0_addr),
    .R0_clk(mem_208_7_R0_clk),
    .R0_data(mem_208_7_R0_data),
    .R0_en(mem_208_7_R0_en),
    .W0_addr(mem_208_7_W0_addr),
    .W0_clk(mem_208_7_W0_clk),
    .W0_data(mem_208_7_W0_data),
    .W0_en(mem_208_7_W0_en),
    .W0_mask(mem_208_7_W0_mask)
  );
  split_mem_0_ext mem_209_0 (
    .R0_addr(mem_209_0_R0_addr),
    .R0_clk(mem_209_0_R0_clk),
    .R0_data(mem_209_0_R0_data),
    .R0_en(mem_209_0_R0_en),
    .W0_addr(mem_209_0_W0_addr),
    .W0_clk(mem_209_0_W0_clk),
    .W0_data(mem_209_0_W0_data),
    .W0_en(mem_209_0_W0_en),
    .W0_mask(mem_209_0_W0_mask)
  );
  split_mem_0_ext mem_209_1 (
    .R0_addr(mem_209_1_R0_addr),
    .R0_clk(mem_209_1_R0_clk),
    .R0_data(mem_209_1_R0_data),
    .R0_en(mem_209_1_R0_en),
    .W0_addr(mem_209_1_W0_addr),
    .W0_clk(mem_209_1_W0_clk),
    .W0_data(mem_209_1_W0_data),
    .W0_en(mem_209_1_W0_en),
    .W0_mask(mem_209_1_W0_mask)
  );
  split_mem_0_ext mem_209_2 (
    .R0_addr(mem_209_2_R0_addr),
    .R0_clk(mem_209_2_R0_clk),
    .R0_data(mem_209_2_R0_data),
    .R0_en(mem_209_2_R0_en),
    .W0_addr(mem_209_2_W0_addr),
    .W0_clk(mem_209_2_W0_clk),
    .W0_data(mem_209_2_W0_data),
    .W0_en(mem_209_2_W0_en),
    .W0_mask(mem_209_2_W0_mask)
  );
  split_mem_0_ext mem_209_3 (
    .R0_addr(mem_209_3_R0_addr),
    .R0_clk(mem_209_3_R0_clk),
    .R0_data(mem_209_3_R0_data),
    .R0_en(mem_209_3_R0_en),
    .W0_addr(mem_209_3_W0_addr),
    .W0_clk(mem_209_3_W0_clk),
    .W0_data(mem_209_3_W0_data),
    .W0_en(mem_209_3_W0_en),
    .W0_mask(mem_209_3_W0_mask)
  );
  split_mem_0_ext mem_209_4 (
    .R0_addr(mem_209_4_R0_addr),
    .R0_clk(mem_209_4_R0_clk),
    .R0_data(mem_209_4_R0_data),
    .R0_en(mem_209_4_R0_en),
    .W0_addr(mem_209_4_W0_addr),
    .W0_clk(mem_209_4_W0_clk),
    .W0_data(mem_209_4_W0_data),
    .W0_en(mem_209_4_W0_en),
    .W0_mask(mem_209_4_W0_mask)
  );
  split_mem_0_ext mem_209_5 (
    .R0_addr(mem_209_5_R0_addr),
    .R0_clk(mem_209_5_R0_clk),
    .R0_data(mem_209_5_R0_data),
    .R0_en(mem_209_5_R0_en),
    .W0_addr(mem_209_5_W0_addr),
    .W0_clk(mem_209_5_W0_clk),
    .W0_data(mem_209_5_W0_data),
    .W0_en(mem_209_5_W0_en),
    .W0_mask(mem_209_5_W0_mask)
  );
  split_mem_0_ext mem_209_6 (
    .R0_addr(mem_209_6_R0_addr),
    .R0_clk(mem_209_6_R0_clk),
    .R0_data(mem_209_6_R0_data),
    .R0_en(mem_209_6_R0_en),
    .W0_addr(mem_209_6_W0_addr),
    .W0_clk(mem_209_6_W0_clk),
    .W0_data(mem_209_6_W0_data),
    .W0_en(mem_209_6_W0_en),
    .W0_mask(mem_209_6_W0_mask)
  );
  split_mem_0_ext mem_209_7 (
    .R0_addr(mem_209_7_R0_addr),
    .R0_clk(mem_209_7_R0_clk),
    .R0_data(mem_209_7_R0_data),
    .R0_en(mem_209_7_R0_en),
    .W0_addr(mem_209_7_W0_addr),
    .W0_clk(mem_209_7_W0_clk),
    .W0_data(mem_209_7_W0_data),
    .W0_en(mem_209_7_W0_en),
    .W0_mask(mem_209_7_W0_mask)
  );
  split_mem_0_ext mem_210_0 (
    .R0_addr(mem_210_0_R0_addr),
    .R0_clk(mem_210_0_R0_clk),
    .R0_data(mem_210_0_R0_data),
    .R0_en(mem_210_0_R0_en),
    .W0_addr(mem_210_0_W0_addr),
    .W0_clk(mem_210_0_W0_clk),
    .W0_data(mem_210_0_W0_data),
    .W0_en(mem_210_0_W0_en),
    .W0_mask(mem_210_0_W0_mask)
  );
  split_mem_0_ext mem_210_1 (
    .R0_addr(mem_210_1_R0_addr),
    .R0_clk(mem_210_1_R0_clk),
    .R0_data(mem_210_1_R0_data),
    .R0_en(mem_210_1_R0_en),
    .W0_addr(mem_210_1_W0_addr),
    .W0_clk(mem_210_1_W0_clk),
    .W0_data(mem_210_1_W0_data),
    .W0_en(mem_210_1_W0_en),
    .W0_mask(mem_210_1_W0_mask)
  );
  split_mem_0_ext mem_210_2 (
    .R0_addr(mem_210_2_R0_addr),
    .R0_clk(mem_210_2_R0_clk),
    .R0_data(mem_210_2_R0_data),
    .R0_en(mem_210_2_R0_en),
    .W0_addr(mem_210_2_W0_addr),
    .W0_clk(mem_210_2_W0_clk),
    .W0_data(mem_210_2_W0_data),
    .W0_en(mem_210_2_W0_en),
    .W0_mask(mem_210_2_W0_mask)
  );
  split_mem_0_ext mem_210_3 (
    .R0_addr(mem_210_3_R0_addr),
    .R0_clk(mem_210_3_R0_clk),
    .R0_data(mem_210_3_R0_data),
    .R0_en(mem_210_3_R0_en),
    .W0_addr(mem_210_3_W0_addr),
    .W0_clk(mem_210_3_W0_clk),
    .W0_data(mem_210_3_W0_data),
    .W0_en(mem_210_3_W0_en),
    .W0_mask(mem_210_3_W0_mask)
  );
  split_mem_0_ext mem_210_4 (
    .R0_addr(mem_210_4_R0_addr),
    .R0_clk(mem_210_4_R0_clk),
    .R0_data(mem_210_4_R0_data),
    .R0_en(mem_210_4_R0_en),
    .W0_addr(mem_210_4_W0_addr),
    .W0_clk(mem_210_4_W0_clk),
    .W0_data(mem_210_4_W0_data),
    .W0_en(mem_210_4_W0_en),
    .W0_mask(mem_210_4_W0_mask)
  );
  split_mem_0_ext mem_210_5 (
    .R0_addr(mem_210_5_R0_addr),
    .R0_clk(mem_210_5_R0_clk),
    .R0_data(mem_210_5_R0_data),
    .R0_en(mem_210_5_R0_en),
    .W0_addr(mem_210_5_W0_addr),
    .W0_clk(mem_210_5_W0_clk),
    .W0_data(mem_210_5_W0_data),
    .W0_en(mem_210_5_W0_en),
    .W0_mask(mem_210_5_W0_mask)
  );
  split_mem_0_ext mem_210_6 (
    .R0_addr(mem_210_6_R0_addr),
    .R0_clk(mem_210_6_R0_clk),
    .R0_data(mem_210_6_R0_data),
    .R0_en(mem_210_6_R0_en),
    .W0_addr(mem_210_6_W0_addr),
    .W0_clk(mem_210_6_W0_clk),
    .W0_data(mem_210_6_W0_data),
    .W0_en(mem_210_6_W0_en),
    .W0_mask(mem_210_6_W0_mask)
  );
  split_mem_0_ext mem_210_7 (
    .R0_addr(mem_210_7_R0_addr),
    .R0_clk(mem_210_7_R0_clk),
    .R0_data(mem_210_7_R0_data),
    .R0_en(mem_210_7_R0_en),
    .W0_addr(mem_210_7_W0_addr),
    .W0_clk(mem_210_7_W0_clk),
    .W0_data(mem_210_7_W0_data),
    .W0_en(mem_210_7_W0_en),
    .W0_mask(mem_210_7_W0_mask)
  );
  split_mem_0_ext mem_211_0 (
    .R0_addr(mem_211_0_R0_addr),
    .R0_clk(mem_211_0_R0_clk),
    .R0_data(mem_211_0_R0_data),
    .R0_en(mem_211_0_R0_en),
    .W0_addr(mem_211_0_W0_addr),
    .W0_clk(mem_211_0_W0_clk),
    .W0_data(mem_211_0_W0_data),
    .W0_en(mem_211_0_W0_en),
    .W0_mask(mem_211_0_W0_mask)
  );
  split_mem_0_ext mem_211_1 (
    .R0_addr(mem_211_1_R0_addr),
    .R0_clk(mem_211_1_R0_clk),
    .R0_data(mem_211_1_R0_data),
    .R0_en(mem_211_1_R0_en),
    .W0_addr(mem_211_1_W0_addr),
    .W0_clk(mem_211_1_W0_clk),
    .W0_data(mem_211_1_W0_data),
    .W0_en(mem_211_1_W0_en),
    .W0_mask(mem_211_1_W0_mask)
  );
  split_mem_0_ext mem_211_2 (
    .R0_addr(mem_211_2_R0_addr),
    .R0_clk(mem_211_2_R0_clk),
    .R0_data(mem_211_2_R0_data),
    .R0_en(mem_211_2_R0_en),
    .W0_addr(mem_211_2_W0_addr),
    .W0_clk(mem_211_2_W0_clk),
    .W0_data(mem_211_2_W0_data),
    .W0_en(mem_211_2_W0_en),
    .W0_mask(mem_211_2_W0_mask)
  );
  split_mem_0_ext mem_211_3 (
    .R0_addr(mem_211_3_R0_addr),
    .R0_clk(mem_211_3_R0_clk),
    .R0_data(mem_211_3_R0_data),
    .R0_en(mem_211_3_R0_en),
    .W0_addr(mem_211_3_W0_addr),
    .W0_clk(mem_211_3_W0_clk),
    .W0_data(mem_211_3_W0_data),
    .W0_en(mem_211_3_W0_en),
    .W0_mask(mem_211_3_W0_mask)
  );
  split_mem_0_ext mem_211_4 (
    .R0_addr(mem_211_4_R0_addr),
    .R0_clk(mem_211_4_R0_clk),
    .R0_data(mem_211_4_R0_data),
    .R0_en(mem_211_4_R0_en),
    .W0_addr(mem_211_4_W0_addr),
    .W0_clk(mem_211_4_W0_clk),
    .W0_data(mem_211_4_W0_data),
    .W0_en(mem_211_4_W0_en),
    .W0_mask(mem_211_4_W0_mask)
  );
  split_mem_0_ext mem_211_5 (
    .R0_addr(mem_211_5_R0_addr),
    .R0_clk(mem_211_5_R0_clk),
    .R0_data(mem_211_5_R0_data),
    .R0_en(mem_211_5_R0_en),
    .W0_addr(mem_211_5_W0_addr),
    .W0_clk(mem_211_5_W0_clk),
    .W0_data(mem_211_5_W0_data),
    .W0_en(mem_211_5_W0_en),
    .W0_mask(mem_211_5_W0_mask)
  );
  split_mem_0_ext mem_211_6 (
    .R0_addr(mem_211_6_R0_addr),
    .R0_clk(mem_211_6_R0_clk),
    .R0_data(mem_211_6_R0_data),
    .R0_en(mem_211_6_R0_en),
    .W0_addr(mem_211_6_W0_addr),
    .W0_clk(mem_211_6_W0_clk),
    .W0_data(mem_211_6_W0_data),
    .W0_en(mem_211_6_W0_en),
    .W0_mask(mem_211_6_W0_mask)
  );
  split_mem_0_ext mem_211_7 (
    .R0_addr(mem_211_7_R0_addr),
    .R0_clk(mem_211_7_R0_clk),
    .R0_data(mem_211_7_R0_data),
    .R0_en(mem_211_7_R0_en),
    .W0_addr(mem_211_7_W0_addr),
    .W0_clk(mem_211_7_W0_clk),
    .W0_data(mem_211_7_W0_data),
    .W0_en(mem_211_7_W0_en),
    .W0_mask(mem_211_7_W0_mask)
  );
  split_mem_0_ext mem_212_0 (
    .R0_addr(mem_212_0_R0_addr),
    .R0_clk(mem_212_0_R0_clk),
    .R0_data(mem_212_0_R0_data),
    .R0_en(mem_212_0_R0_en),
    .W0_addr(mem_212_0_W0_addr),
    .W0_clk(mem_212_0_W0_clk),
    .W0_data(mem_212_0_W0_data),
    .W0_en(mem_212_0_W0_en),
    .W0_mask(mem_212_0_W0_mask)
  );
  split_mem_0_ext mem_212_1 (
    .R0_addr(mem_212_1_R0_addr),
    .R0_clk(mem_212_1_R0_clk),
    .R0_data(mem_212_1_R0_data),
    .R0_en(mem_212_1_R0_en),
    .W0_addr(mem_212_1_W0_addr),
    .W0_clk(mem_212_1_W0_clk),
    .W0_data(mem_212_1_W0_data),
    .W0_en(mem_212_1_W0_en),
    .W0_mask(mem_212_1_W0_mask)
  );
  split_mem_0_ext mem_212_2 (
    .R0_addr(mem_212_2_R0_addr),
    .R0_clk(mem_212_2_R0_clk),
    .R0_data(mem_212_2_R0_data),
    .R0_en(mem_212_2_R0_en),
    .W0_addr(mem_212_2_W0_addr),
    .W0_clk(mem_212_2_W0_clk),
    .W0_data(mem_212_2_W0_data),
    .W0_en(mem_212_2_W0_en),
    .W0_mask(mem_212_2_W0_mask)
  );
  split_mem_0_ext mem_212_3 (
    .R0_addr(mem_212_3_R0_addr),
    .R0_clk(mem_212_3_R0_clk),
    .R0_data(mem_212_3_R0_data),
    .R0_en(mem_212_3_R0_en),
    .W0_addr(mem_212_3_W0_addr),
    .W0_clk(mem_212_3_W0_clk),
    .W0_data(mem_212_3_W0_data),
    .W0_en(mem_212_3_W0_en),
    .W0_mask(mem_212_3_W0_mask)
  );
  split_mem_0_ext mem_212_4 (
    .R0_addr(mem_212_4_R0_addr),
    .R0_clk(mem_212_4_R0_clk),
    .R0_data(mem_212_4_R0_data),
    .R0_en(mem_212_4_R0_en),
    .W0_addr(mem_212_4_W0_addr),
    .W0_clk(mem_212_4_W0_clk),
    .W0_data(mem_212_4_W0_data),
    .W0_en(mem_212_4_W0_en),
    .W0_mask(mem_212_4_W0_mask)
  );
  split_mem_0_ext mem_212_5 (
    .R0_addr(mem_212_5_R0_addr),
    .R0_clk(mem_212_5_R0_clk),
    .R0_data(mem_212_5_R0_data),
    .R0_en(mem_212_5_R0_en),
    .W0_addr(mem_212_5_W0_addr),
    .W0_clk(mem_212_5_W0_clk),
    .W0_data(mem_212_5_W0_data),
    .W0_en(mem_212_5_W0_en),
    .W0_mask(mem_212_5_W0_mask)
  );
  split_mem_0_ext mem_212_6 (
    .R0_addr(mem_212_6_R0_addr),
    .R0_clk(mem_212_6_R0_clk),
    .R0_data(mem_212_6_R0_data),
    .R0_en(mem_212_6_R0_en),
    .W0_addr(mem_212_6_W0_addr),
    .W0_clk(mem_212_6_W0_clk),
    .W0_data(mem_212_6_W0_data),
    .W0_en(mem_212_6_W0_en),
    .W0_mask(mem_212_6_W0_mask)
  );
  split_mem_0_ext mem_212_7 (
    .R0_addr(mem_212_7_R0_addr),
    .R0_clk(mem_212_7_R0_clk),
    .R0_data(mem_212_7_R0_data),
    .R0_en(mem_212_7_R0_en),
    .W0_addr(mem_212_7_W0_addr),
    .W0_clk(mem_212_7_W0_clk),
    .W0_data(mem_212_7_W0_data),
    .W0_en(mem_212_7_W0_en),
    .W0_mask(mem_212_7_W0_mask)
  );
  split_mem_0_ext mem_213_0 (
    .R0_addr(mem_213_0_R0_addr),
    .R0_clk(mem_213_0_R0_clk),
    .R0_data(mem_213_0_R0_data),
    .R0_en(mem_213_0_R0_en),
    .W0_addr(mem_213_0_W0_addr),
    .W0_clk(mem_213_0_W0_clk),
    .W0_data(mem_213_0_W0_data),
    .W0_en(mem_213_0_W0_en),
    .W0_mask(mem_213_0_W0_mask)
  );
  split_mem_0_ext mem_213_1 (
    .R0_addr(mem_213_1_R0_addr),
    .R0_clk(mem_213_1_R0_clk),
    .R0_data(mem_213_1_R0_data),
    .R0_en(mem_213_1_R0_en),
    .W0_addr(mem_213_1_W0_addr),
    .W0_clk(mem_213_1_W0_clk),
    .W0_data(mem_213_1_W0_data),
    .W0_en(mem_213_1_W0_en),
    .W0_mask(mem_213_1_W0_mask)
  );
  split_mem_0_ext mem_213_2 (
    .R0_addr(mem_213_2_R0_addr),
    .R0_clk(mem_213_2_R0_clk),
    .R0_data(mem_213_2_R0_data),
    .R0_en(mem_213_2_R0_en),
    .W0_addr(mem_213_2_W0_addr),
    .W0_clk(mem_213_2_W0_clk),
    .W0_data(mem_213_2_W0_data),
    .W0_en(mem_213_2_W0_en),
    .W0_mask(mem_213_2_W0_mask)
  );
  split_mem_0_ext mem_213_3 (
    .R0_addr(mem_213_3_R0_addr),
    .R0_clk(mem_213_3_R0_clk),
    .R0_data(mem_213_3_R0_data),
    .R0_en(mem_213_3_R0_en),
    .W0_addr(mem_213_3_W0_addr),
    .W0_clk(mem_213_3_W0_clk),
    .W0_data(mem_213_3_W0_data),
    .W0_en(mem_213_3_W0_en),
    .W0_mask(mem_213_3_W0_mask)
  );
  split_mem_0_ext mem_213_4 (
    .R0_addr(mem_213_4_R0_addr),
    .R0_clk(mem_213_4_R0_clk),
    .R0_data(mem_213_4_R0_data),
    .R0_en(mem_213_4_R0_en),
    .W0_addr(mem_213_4_W0_addr),
    .W0_clk(mem_213_4_W0_clk),
    .W0_data(mem_213_4_W0_data),
    .W0_en(mem_213_4_W0_en),
    .W0_mask(mem_213_4_W0_mask)
  );
  split_mem_0_ext mem_213_5 (
    .R0_addr(mem_213_5_R0_addr),
    .R0_clk(mem_213_5_R0_clk),
    .R0_data(mem_213_5_R0_data),
    .R0_en(mem_213_5_R0_en),
    .W0_addr(mem_213_5_W0_addr),
    .W0_clk(mem_213_5_W0_clk),
    .W0_data(mem_213_5_W0_data),
    .W0_en(mem_213_5_W0_en),
    .W0_mask(mem_213_5_W0_mask)
  );
  split_mem_0_ext mem_213_6 (
    .R0_addr(mem_213_6_R0_addr),
    .R0_clk(mem_213_6_R0_clk),
    .R0_data(mem_213_6_R0_data),
    .R0_en(mem_213_6_R0_en),
    .W0_addr(mem_213_6_W0_addr),
    .W0_clk(mem_213_6_W0_clk),
    .W0_data(mem_213_6_W0_data),
    .W0_en(mem_213_6_W0_en),
    .W0_mask(mem_213_6_W0_mask)
  );
  split_mem_0_ext mem_213_7 (
    .R0_addr(mem_213_7_R0_addr),
    .R0_clk(mem_213_7_R0_clk),
    .R0_data(mem_213_7_R0_data),
    .R0_en(mem_213_7_R0_en),
    .W0_addr(mem_213_7_W0_addr),
    .W0_clk(mem_213_7_W0_clk),
    .W0_data(mem_213_7_W0_data),
    .W0_en(mem_213_7_W0_en),
    .W0_mask(mem_213_7_W0_mask)
  );
  split_mem_0_ext mem_214_0 (
    .R0_addr(mem_214_0_R0_addr),
    .R0_clk(mem_214_0_R0_clk),
    .R0_data(mem_214_0_R0_data),
    .R0_en(mem_214_0_R0_en),
    .W0_addr(mem_214_0_W0_addr),
    .W0_clk(mem_214_0_W0_clk),
    .W0_data(mem_214_0_W0_data),
    .W0_en(mem_214_0_W0_en),
    .W0_mask(mem_214_0_W0_mask)
  );
  split_mem_0_ext mem_214_1 (
    .R0_addr(mem_214_1_R0_addr),
    .R0_clk(mem_214_1_R0_clk),
    .R0_data(mem_214_1_R0_data),
    .R0_en(mem_214_1_R0_en),
    .W0_addr(mem_214_1_W0_addr),
    .W0_clk(mem_214_1_W0_clk),
    .W0_data(mem_214_1_W0_data),
    .W0_en(mem_214_1_W0_en),
    .W0_mask(mem_214_1_W0_mask)
  );
  split_mem_0_ext mem_214_2 (
    .R0_addr(mem_214_2_R0_addr),
    .R0_clk(mem_214_2_R0_clk),
    .R0_data(mem_214_2_R0_data),
    .R0_en(mem_214_2_R0_en),
    .W0_addr(mem_214_2_W0_addr),
    .W0_clk(mem_214_2_W0_clk),
    .W0_data(mem_214_2_W0_data),
    .W0_en(mem_214_2_W0_en),
    .W0_mask(mem_214_2_W0_mask)
  );
  split_mem_0_ext mem_214_3 (
    .R0_addr(mem_214_3_R0_addr),
    .R0_clk(mem_214_3_R0_clk),
    .R0_data(mem_214_3_R0_data),
    .R0_en(mem_214_3_R0_en),
    .W0_addr(mem_214_3_W0_addr),
    .W0_clk(mem_214_3_W0_clk),
    .W0_data(mem_214_3_W0_data),
    .W0_en(mem_214_3_W0_en),
    .W0_mask(mem_214_3_W0_mask)
  );
  split_mem_0_ext mem_214_4 (
    .R0_addr(mem_214_4_R0_addr),
    .R0_clk(mem_214_4_R0_clk),
    .R0_data(mem_214_4_R0_data),
    .R0_en(mem_214_4_R0_en),
    .W0_addr(mem_214_4_W0_addr),
    .W0_clk(mem_214_4_W0_clk),
    .W0_data(mem_214_4_W0_data),
    .W0_en(mem_214_4_W0_en),
    .W0_mask(mem_214_4_W0_mask)
  );
  split_mem_0_ext mem_214_5 (
    .R0_addr(mem_214_5_R0_addr),
    .R0_clk(mem_214_5_R0_clk),
    .R0_data(mem_214_5_R0_data),
    .R0_en(mem_214_5_R0_en),
    .W0_addr(mem_214_5_W0_addr),
    .W0_clk(mem_214_5_W0_clk),
    .W0_data(mem_214_5_W0_data),
    .W0_en(mem_214_5_W0_en),
    .W0_mask(mem_214_5_W0_mask)
  );
  split_mem_0_ext mem_214_6 (
    .R0_addr(mem_214_6_R0_addr),
    .R0_clk(mem_214_6_R0_clk),
    .R0_data(mem_214_6_R0_data),
    .R0_en(mem_214_6_R0_en),
    .W0_addr(mem_214_6_W0_addr),
    .W0_clk(mem_214_6_W0_clk),
    .W0_data(mem_214_6_W0_data),
    .W0_en(mem_214_6_W0_en),
    .W0_mask(mem_214_6_W0_mask)
  );
  split_mem_0_ext mem_214_7 (
    .R0_addr(mem_214_7_R0_addr),
    .R0_clk(mem_214_7_R0_clk),
    .R0_data(mem_214_7_R0_data),
    .R0_en(mem_214_7_R0_en),
    .W0_addr(mem_214_7_W0_addr),
    .W0_clk(mem_214_7_W0_clk),
    .W0_data(mem_214_7_W0_data),
    .W0_en(mem_214_7_W0_en),
    .W0_mask(mem_214_7_W0_mask)
  );
  split_mem_0_ext mem_215_0 (
    .R0_addr(mem_215_0_R0_addr),
    .R0_clk(mem_215_0_R0_clk),
    .R0_data(mem_215_0_R0_data),
    .R0_en(mem_215_0_R0_en),
    .W0_addr(mem_215_0_W0_addr),
    .W0_clk(mem_215_0_W0_clk),
    .W0_data(mem_215_0_W0_data),
    .W0_en(mem_215_0_W0_en),
    .W0_mask(mem_215_0_W0_mask)
  );
  split_mem_0_ext mem_215_1 (
    .R0_addr(mem_215_1_R0_addr),
    .R0_clk(mem_215_1_R0_clk),
    .R0_data(mem_215_1_R0_data),
    .R0_en(mem_215_1_R0_en),
    .W0_addr(mem_215_1_W0_addr),
    .W0_clk(mem_215_1_W0_clk),
    .W0_data(mem_215_1_W0_data),
    .W0_en(mem_215_1_W0_en),
    .W0_mask(mem_215_1_W0_mask)
  );
  split_mem_0_ext mem_215_2 (
    .R0_addr(mem_215_2_R0_addr),
    .R0_clk(mem_215_2_R0_clk),
    .R0_data(mem_215_2_R0_data),
    .R0_en(mem_215_2_R0_en),
    .W0_addr(mem_215_2_W0_addr),
    .W0_clk(mem_215_2_W0_clk),
    .W0_data(mem_215_2_W0_data),
    .W0_en(mem_215_2_W0_en),
    .W0_mask(mem_215_2_W0_mask)
  );
  split_mem_0_ext mem_215_3 (
    .R0_addr(mem_215_3_R0_addr),
    .R0_clk(mem_215_3_R0_clk),
    .R0_data(mem_215_3_R0_data),
    .R0_en(mem_215_3_R0_en),
    .W0_addr(mem_215_3_W0_addr),
    .W0_clk(mem_215_3_W0_clk),
    .W0_data(mem_215_3_W0_data),
    .W0_en(mem_215_3_W0_en),
    .W0_mask(mem_215_3_W0_mask)
  );
  split_mem_0_ext mem_215_4 (
    .R0_addr(mem_215_4_R0_addr),
    .R0_clk(mem_215_4_R0_clk),
    .R0_data(mem_215_4_R0_data),
    .R0_en(mem_215_4_R0_en),
    .W0_addr(mem_215_4_W0_addr),
    .W0_clk(mem_215_4_W0_clk),
    .W0_data(mem_215_4_W0_data),
    .W0_en(mem_215_4_W0_en),
    .W0_mask(mem_215_4_W0_mask)
  );
  split_mem_0_ext mem_215_5 (
    .R0_addr(mem_215_5_R0_addr),
    .R0_clk(mem_215_5_R0_clk),
    .R0_data(mem_215_5_R0_data),
    .R0_en(mem_215_5_R0_en),
    .W0_addr(mem_215_5_W0_addr),
    .W0_clk(mem_215_5_W0_clk),
    .W0_data(mem_215_5_W0_data),
    .W0_en(mem_215_5_W0_en),
    .W0_mask(mem_215_5_W0_mask)
  );
  split_mem_0_ext mem_215_6 (
    .R0_addr(mem_215_6_R0_addr),
    .R0_clk(mem_215_6_R0_clk),
    .R0_data(mem_215_6_R0_data),
    .R0_en(mem_215_6_R0_en),
    .W0_addr(mem_215_6_W0_addr),
    .W0_clk(mem_215_6_W0_clk),
    .W0_data(mem_215_6_W0_data),
    .W0_en(mem_215_6_W0_en),
    .W0_mask(mem_215_6_W0_mask)
  );
  split_mem_0_ext mem_215_7 (
    .R0_addr(mem_215_7_R0_addr),
    .R0_clk(mem_215_7_R0_clk),
    .R0_data(mem_215_7_R0_data),
    .R0_en(mem_215_7_R0_en),
    .W0_addr(mem_215_7_W0_addr),
    .W0_clk(mem_215_7_W0_clk),
    .W0_data(mem_215_7_W0_data),
    .W0_en(mem_215_7_W0_en),
    .W0_mask(mem_215_7_W0_mask)
  );
  split_mem_0_ext mem_216_0 (
    .R0_addr(mem_216_0_R0_addr),
    .R0_clk(mem_216_0_R0_clk),
    .R0_data(mem_216_0_R0_data),
    .R0_en(mem_216_0_R0_en),
    .W0_addr(mem_216_0_W0_addr),
    .W0_clk(mem_216_0_W0_clk),
    .W0_data(mem_216_0_W0_data),
    .W0_en(mem_216_0_W0_en),
    .W0_mask(mem_216_0_W0_mask)
  );
  split_mem_0_ext mem_216_1 (
    .R0_addr(mem_216_1_R0_addr),
    .R0_clk(mem_216_1_R0_clk),
    .R0_data(mem_216_1_R0_data),
    .R0_en(mem_216_1_R0_en),
    .W0_addr(mem_216_1_W0_addr),
    .W0_clk(mem_216_1_W0_clk),
    .W0_data(mem_216_1_W0_data),
    .W0_en(mem_216_1_W0_en),
    .W0_mask(mem_216_1_W0_mask)
  );
  split_mem_0_ext mem_216_2 (
    .R0_addr(mem_216_2_R0_addr),
    .R0_clk(mem_216_2_R0_clk),
    .R0_data(mem_216_2_R0_data),
    .R0_en(mem_216_2_R0_en),
    .W0_addr(mem_216_2_W0_addr),
    .W0_clk(mem_216_2_W0_clk),
    .W0_data(mem_216_2_W0_data),
    .W0_en(mem_216_2_W0_en),
    .W0_mask(mem_216_2_W0_mask)
  );
  split_mem_0_ext mem_216_3 (
    .R0_addr(mem_216_3_R0_addr),
    .R0_clk(mem_216_3_R0_clk),
    .R0_data(mem_216_3_R0_data),
    .R0_en(mem_216_3_R0_en),
    .W0_addr(mem_216_3_W0_addr),
    .W0_clk(mem_216_3_W0_clk),
    .W0_data(mem_216_3_W0_data),
    .W0_en(mem_216_3_W0_en),
    .W0_mask(mem_216_3_W0_mask)
  );
  split_mem_0_ext mem_216_4 (
    .R0_addr(mem_216_4_R0_addr),
    .R0_clk(mem_216_4_R0_clk),
    .R0_data(mem_216_4_R0_data),
    .R0_en(mem_216_4_R0_en),
    .W0_addr(mem_216_4_W0_addr),
    .W0_clk(mem_216_4_W0_clk),
    .W0_data(mem_216_4_W0_data),
    .W0_en(mem_216_4_W0_en),
    .W0_mask(mem_216_4_W0_mask)
  );
  split_mem_0_ext mem_216_5 (
    .R0_addr(mem_216_5_R0_addr),
    .R0_clk(mem_216_5_R0_clk),
    .R0_data(mem_216_5_R0_data),
    .R0_en(mem_216_5_R0_en),
    .W0_addr(mem_216_5_W0_addr),
    .W0_clk(mem_216_5_W0_clk),
    .W0_data(mem_216_5_W0_data),
    .W0_en(mem_216_5_W0_en),
    .W0_mask(mem_216_5_W0_mask)
  );
  split_mem_0_ext mem_216_6 (
    .R0_addr(mem_216_6_R0_addr),
    .R0_clk(mem_216_6_R0_clk),
    .R0_data(mem_216_6_R0_data),
    .R0_en(mem_216_6_R0_en),
    .W0_addr(mem_216_6_W0_addr),
    .W0_clk(mem_216_6_W0_clk),
    .W0_data(mem_216_6_W0_data),
    .W0_en(mem_216_6_W0_en),
    .W0_mask(mem_216_6_W0_mask)
  );
  split_mem_0_ext mem_216_7 (
    .R0_addr(mem_216_7_R0_addr),
    .R0_clk(mem_216_7_R0_clk),
    .R0_data(mem_216_7_R0_data),
    .R0_en(mem_216_7_R0_en),
    .W0_addr(mem_216_7_W0_addr),
    .W0_clk(mem_216_7_W0_clk),
    .W0_data(mem_216_7_W0_data),
    .W0_en(mem_216_7_W0_en),
    .W0_mask(mem_216_7_W0_mask)
  );
  split_mem_0_ext mem_217_0 (
    .R0_addr(mem_217_0_R0_addr),
    .R0_clk(mem_217_0_R0_clk),
    .R0_data(mem_217_0_R0_data),
    .R0_en(mem_217_0_R0_en),
    .W0_addr(mem_217_0_W0_addr),
    .W0_clk(mem_217_0_W0_clk),
    .W0_data(mem_217_0_W0_data),
    .W0_en(mem_217_0_W0_en),
    .W0_mask(mem_217_0_W0_mask)
  );
  split_mem_0_ext mem_217_1 (
    .R0_addr(mem_217_1_R0_addr),
    .R0_clk(mem_217_1_R0_clk),
    .R0_data(mem_217_1_R0_data),
    .R0_en(mem_217_1_R0_en),
    .W0_addr(mem_217_1_W0_addr),
    .W0_clk(mem_217_1_W0_clk),
    .W0_data(mem_217_1_W0_data),
    .W0_en(mem_217_1_W0_en),
    .W0_mask(mem_217_1_W0_mask)
  );
  split_mem_0_ext mem_217_2 (
    .R0_addr(mem_217_2_R0_addr),
    .R0_clk(mem_217_2_R0_clk),
    .R0_data(mem_217_2_R0_data),
    .R0_en(mem_217_2_R0_en),
    .W0_addr(mem_217_2_W0_addr),
    .W0_clk(mem_217_2_W0_clk),
    .W0_data(mem_217_2_W0_data),
    .W0_en(mem_217_2_W0_en),
    .W0_mask(mem_217_2_W0_mask)
  );
  split_mem_0_ext mem_217_3 (
    .R0_addr(mem_217_3_R0_addr),
    .R0_clk(mem_217_3_R0_clk),
    .R0_data(mem_217_3_R0_data),
    .R0_en(mem_217_3_R0_en),
    .W0_addr(mem_217_3_W0_addr),
    .W0_clk(mem_217_3_W0_clk),
    .W0_data(mem_217_3_W0_data),
    .W0_en(mem_217_3_W0_en),
    .W0_mask(mem_217_3_W0_mask)
  );
  split_mem_0_ext mem_217_4 (
    .R0_addr(mem_217_4_R0_addr),
    .R0_clk(mem_217_4_R0_clk),
    .R0_data(mem_217_4_R0_data),
    .R0_en(mem_217_4_R0_en),
    .W0_addr(mem_217_4_W0_addr),
    .W0_clk(mem_217_4_W0_clk),
    .W0_data(mem_217_4_W0_data),
    .W0_en(mem_217_4_W0_en),
    .W0_mask(mem_217_4_W0_mask)
  );
  split_mem_0_ext mem_217_5 (
    .R0_addr(mem_217_5_R0_addr),
    .R0_clk(mem_217_5_R0_clk),
    .R0_data(mem_217_5_R0_data),
    .R0_en(mem_217_5_R0_en),
    .W0_addr(mem_217_5_W0_addr),
    .W0_clk(mem_217_5_W0_clk),
    .W0_data(mem_217_5_W0_data),
    .W0_en(mem_217_5_W0_en),
    .W0_mask(mem_217_5_W0_mask)
  );
  split_mem_0_ext mem_217_6 (
    .R0_addr(mem_217_6_R0_addr),
    .R0_clk(mem_217_6_R0_clk),
    .R0_data(mem_217_6_R0_data),
    .R0_en(mem_217_6_R0_en),
    .W0_addr(mem_217_6_W0_addr),
    .W0_clk(mem_217_6_W0_clk),
    .W0_data(mem_217_6_W0_data),
    .W0_en(mem_217_6_W0_en),
    .W0_mask(mem_217_6_W0_mask)
  );
  split_mem_0_ext mem_217_7 (
    .R0_addr(mem_217_7_R0_addr),
    .R0_clk(mem_217_7_R0_clk),
    .R0_data(mem_217_7_R0_data),
    .R0_en(mem_217_7_R0_en),
    .W0_addr(mem_217_7_W0_addr),
    .W0_clk(mem_217_7_W0_clk),
    .W0_data(mem_217_7_W0_data),
    .W0_en(mem_217_7_W0_en),
    .W0_mask(mem_217_7_W0_mask)
  );
  split_mem_0_ext mem_218_0 (
    .R0_addr(mem_218_0_R0_addr),
    .R0_clk(mem_218_0_R0_clk),
    .R0_data(mem_218_0_R0_data),
    .R0_en(mem_218_0_R0_en),
    .W0_addr(mem_218_0_W0_addr),
    .W0_clk(mem_218_0_W0_clk),
    .W0_data(mem_218_0_W0_data),
    .W0_en(mem_218_0_W0_en),
    .W0_mask(mem_218_0_W0_mask)
  );
  split_mem_0_ext mem_218_1 (
    .R0_addr(mem_218_1_R0_addr),
    .R0_clk(mem_218_1_R0_clk),
    .R0_data(mem_218_1_R0_data),
    .R0_en(mem_218_1_R0_en),
    .W0_addr(mem_218_1_W0_addr),
    .W0_clk(mem_218_1_W0_clk),
    .W0_data(mem_218_1_W0_data),
    .W0_en(mem_218_1_W0_en),
    .W0_mask(mem_218_1_W0_mask)
  );
  split_mem_0_ext mem_218_2 (
    .R0_addr(mem_218_2_R0_addr),
    .R0_clk(mem_218_2_R0_clk),
    .R0_data(mem_218_2_R0_data),
    .R0_en(mem_218_2_R0_en),
    .W0_addr(mem_218_2_W0_addr),
    .W0_clk(mem_218_2_W0_clk),
    .W0_data(mem_218_2_W0_data),
    .W0_en(mem_218_2_W0_en),
    .W0_mask(mem_218_2_W0_mask)
  );
  split_mem_0_ext mem_218_3 (
    .R0_addr(mem_218_3_R0_addr),
    .R0_clk(mem_218_3_R0_clk),
    .R0_data(mem_218_3_R0_data),
    .R0_en(mem_218_3_R0_en),
    .W0_addr(mem_218_3_W0_addr),
    .W0_clk(mem_218_3_W0_clk),
    .W0_data(mem_218_3_W0_data),
    .W0_en(mem_218_3_W0_en),
    .W0_mask(mem_218_3_W0_mask)
  );
  split_mem_0_ext mem_218_4 (
    .R0_addr(mem_218_4_R0_addr),
    .R0_clk(mem_218_4_R0_clk),
    .R0_data(mem_218_4_R0_data),
    .R0_en(mem_218_4_R0_en),
    .W0_addr(mem_218_4_W0_addr),
    .W0_clk(mem_218_4_W0_clk),
    .W0_data(mem_218_4_W0_data),
    .W0_en(mem_218_4_W0_en),
    .W0_mask(mem_218_4_W0_mask)
  );
  split_mem_0_ext mem_218_5 (
    .R0_addr(mem_218_5_R0_addr),
    .R0_clk(mem_218_5_R0_clk),
    .R0_data(mem_218_5_R0_data),
    .R0_en(mem_218_5_R0_en),
    .W0_addr(mem_218_5_W0_addr),
    .W0_clk(mem_218_5_W0_clk),
    .W0_data(mem_218_5_W0_data),
    .W0_en(mem_218_5_W0_en),
    .W0_mask(mem_218_5_W0_mask)
  );
  split_mem_0_ext mem_218_6 (
    .R0_addr(mem_218_6_R0_addr),
    .R0_clk(mem_218_6_R0_clk),
    .R0_data(mem_218_6_R0_data),
    .R0_en(mem_218_6_R0_en),
    .W0_addr(mem_218_6_W0_addr),
    .W0_clk(mem_218_6_W0_clk),
    .W0_data(mem_218_6_W0_data),
    .W0_en(mem_218_6_W0_en),
    .W0_mask(mem_218_6_W0_mask)
  );
  split_mem_0_ext mem_218_7 (
    .R0_addr(mem_218_7_R0_addr),
    .R0_clk(mem_218_7_R0_clk),
    .R0_data(mem_218_7_R0_data),
    .R0_en(mem_218_7_R0_en),
    .W0_addr(mem_218_7_W0_addr),
    .W0_clk(mem_218_7_W0_clk),
    .W0_data(mem_218_7_W0_data),
    .W0_en(mem_218_7_W0_en),
    .W0_mask(mem_218_7_W0_mask)
  );
  split_mem_0_ext mem_219_0 (
    .R0_addr(mem_219_0_R0_addr),
    .R0_clk(mem_219_0_R0_clk),
    .R0_data(mem_219_0_R0_data),
    .R0_en(mem_219_0_R0_en),
    .W0_addr(mem_219_0_W0_addr),
    .W0_clk(mem_219_0_W0_clk),
    .W0_data(mem_219_0_W0_data),
    .W0_en(mem_219_0_W0_en),
    .W0_mask(mem_219_0_W0_mask)
  );
  split_mem_0_ext mem_219_1 (
    .R0_addr(mem_219_1_R0_addr),
    .R0_clk(mem_219_1_R0_clk),
    .R0_data(mem_219_1_R0_data),
    .R0_en(mem_219_1_R0_en),
    .W0_addr(mem_219_1_W0_addr),
    .W0_clk(mem_219_1_W0_clk),
    .W0_data(mem_219_1_W0_data),
    .W0_en(mem_219_1_W0_en),
    .W0_mask(mem_219_1_W0_mask)
  );
  split_mem_0_ext mem_219_2 (
    .R0_addr(mem_219_2_R0_addr),
    .R0_clk(mem_219_2_R0_clk),
    .R0_data(mem_219_2_R0_data),
    .R0_en(mem_219_2_R0_en),
    .W0_addr(mem_219_2_W0_addr),
    .W0_clk(mem_219_2_W0_clk),
    .W0_data(mem_219_2_W0_data),
    .W0_en(mem_219_2_W0_en),
    .W0_mask(mem_219_2_W0_mask)
  );
  split_mem_0_ext mem_219_3 (
    .R0_addr(mem_219_3_R0_addr),
    .R0_clk(mem_219_3_R0_clk),
    .R0_data(mem_219_3_R0_data),
    .R0_en(mem_219_3_R0_en),
    .W0_addr(mem_219_3_W0_addr),
    .W0_clk(mem_219_3_W0_clk),
    .W0_data(mem_219_3_W0_data),
    .W0_en(mem_219_3_W0_en),
    .W0_mask(mem_219_3_W0_mask)
  );
  split_mem_0_ext mem_219_4 (
    .R0_addr(mem_219_4_R0_addr),
    .R0_clk(mem_219_4_R0_clk),
    .R0_data(mem_219_4_R0_data),
    .R0_en(mem_219_4_R0_en),
    .W0_addr(mem_219_4_W0_addr),
    .W0_clk(mem_219_4_W0_clk),
    .W0_data(mem_219_4_W0_data),
    .W0_en(mem_219_4_W0_en),
    .W0_mask(mem_219_4_W0_mask)
  );
  split_mem_0_ext mem_219_5 (
    .R0_addr(mem_219_5_R0_addr),
    .R0_clk(mem_219_5_R0_clk),
    .R0_data(mem_219_5_R0_data),
    .R0_en(mem_219_5_R0_en),
    .W0_addr(mem_219_5_W0_addr),
    .W0_clk(mem_219_5_W0_clk),
    .W0_data(mem_219_5_W0_data),
    .W0_en(mem_219_5_W0_en),
    .W0_mask(mem_219_5_W0_mask)
  );
  split_mem_0_ext mem_219_6 (
    .R0_addr(mem_219_6_R0_addr),
    .R0_clk(mem_219_6_R0_clk),
    .R0_data(mem_219_6_R0_data),
    .R0_en(mem_219_6_R0_en),
    .W0_addr(mem_219_6_W0_addr),
    .W0_clk(mem_219_6_W0_clk),
    .W0_data(mem_219_6_W0_data),
    .W0_en(mem_219_6_W0_en),
    .W0_mask(mem_219_6_W0_mask)
  );
  split_mem_0_ext mem_219_7 (
    .R0_addr(mem_219_7_R0_addr),
    .R0_clk(mem_219_7_R0_clk),
    .R0_data(mem_219_7_R0_data),
    .R0_en(mem_219_7_R0_en),
    .W0_addr(mem_219_7_W0_addr),
    .W0_clk(mem_219_7_W0_clk),
    .W0_data(mem_219_7_W0_data),
    .W0_en(mem_219_7_W0_en),
    .W0_mask(mem_219_7_W0_mask)
  );
  split_mem_0_ext mem_220_0 (
    .R0_addr(mem_220_0_R0_addr),
    .R0_clk(mem_220_0_R0_clk),
    .R0_data(mem_220_0_R0_data),
    .R0_en(mem_220_0_R0_en),
    .W0_addr(mem_220_0_W0_addr),
    .W0_clk(mem_220_0_W0_clk),
    .W0_data(mem_220_0_W0_data),
    .W0_en(mem_220_0_W0_en),
    .W0_mask(mem_220_0_W0_mask)
  );
  split_mem_0_ext mem_220_1 (
    .R0_addr(mem_220_1_R0_addr),
    .R0_clk(mem_220_1_R0_clk),
    .R0_data(mem_220_1_R0_data),
    .R0_en(mem_220_1_R0_en),
    .W0_addr(mem_220_1_W0_addr),
    .W0_clk(mem_220_1_W0_clk),
    .W0_data(mem_220_1_W0_data),
    .W0_en(mem_220_1_W0_en),
    .W0_mask(mem_220_1_W0_mask)
  );
  split_mem_0_ext mem_220_2 (
    .R0_addr(mem_220_2_R0_addr),
    .R0_clk(mem_220_2_R0_clk),
    .R0_data(mem_220_2_R0_data),
    .R0_en(mem_220_2_R0_en),
    .W0_addr(mem_220_2_W0_addr),
    .W0_clk(mem_220_2_W0_clk),
    .W0_data(mem_220_2_W0_data),
    .W0_en(mem_220_2_W0_en),
    .W0_mask(mem_220_2_W0_mask)
  );
  split_mem_0_ext mem_220_3 (
    .R0_addr(mem_220_3_R0_addr),
    .R0_clk(mem_220_3_R0_clk),
    .R0_data(mem_220_3_R0_data),
    .R0_en(mem_220_3_R0_en),
    .W0_addr(mem_220_3_W0_addr),
    .W0_clk(mem_220_3_W0_clk),
    .W0_data(mem_220_3_W0_data),
    .W0_en(mem_220_3_W0_en),
    .W0_mask(mem_220_3_W0_mask)
  );
  split_mem_0_ext mem_220_4 (
    .R0_addr(mem_220_4_R0_addr),
    .R0_clk(mem_220_4_R0_clk),
    .R0_data(mem_220_4_R0_data),
    .R0_en(mem_220_4_R0_en),
    .W0_addr(mem_220_4_W0_addr),
    .W0_clk(mem_220_4_W0_clk),
    .W0_data(mem_220_4_W0_data),
    .W0_en(mem_220_4_W0_en),
    .W0_mask(mem_220_4_W0_mask)
  );
  split_mem_0_ext mem_220_5 (
    .R0_addr(mem_220_5_R0_addr),
    .R0_clk(mem_220_5_R0_clk),
    .R0_data(mem_220_5_R0_data),
    .R0_en(mem_220_5_R0_en),
    .W0_addr(mem_220_5_W0_addr),
    .W0_clk(mem_220_5_W0_clk),
    .W0_data(mem_220_5_W0_data),
    .W0_en(mem_220_5_W0_en),
    .W0_mask(mem_220_5_W0_mask)
  );
  split_mem_0_ext mem_220_6 (
    .R0_addr(mem_220_6_R0_addr),
    .R0_clk(mem_220_6_R0_clk),
    .R0_data(mem_220_6_R0_data),
    .R0_en(mem_220_6_R0_en),
    .W0_addr(mem_220_6_W0_addr),
    .W0_clk(mem_220_6_W0_clk),
    .W0_data(mem_220_6_W0_data),
    .W0_en(mem_220_6_W0_en),
    .W0_mask(mem_220_6_W0_mask)
  );
  split_mem_0_ext mem_220_7 (
    .R0_addr(mem_220_7_R0_addr),
    .R0_clk(mem_220_7_R0_clk),
    .R0_data(mem_220_7_R0_data),
    .R0_en(mem_220_7_R0_en),
    .W0_addr(mem_220_7_W0_addr),
    .W0_clk(mem_220_7_W0_clk),
    .W0_data(mem_220_7_W0_data),
    .W0_en(mem_220_7_W0_en),
    .W0_mask(mem_220_7_W0_mask)
  );
  split_mem_0_ext mem_221_0 (
    .R0_addr(mem_221_0_R0_addr),
    .R0_clk(mem_221_0_R0_clk),
    .R0_data(mem_221_0_R0_data),
    .R0_en(mem_221_0_R0_en),
    .W0_addr(mem_221_0_W0_addr),
    .W0_clk(mem_221_0_W0_clk),
    .W0_data(mem_221_0_W0_data),
    .W0_en(mem_221_0_W0_en),
    .W0_mask(mem_221_0_W0_mask)
  );
  split_mem_0_ext mem_221_1 (
    .R0_addr(mem_221_1_R0_addr),
    .R0_clk(mem_221_1_R0_clk),
    .R0_data(mem_221_1_R0_data),
    .R0_en(mem_221_1_R0_en),
    .W0_addr(mem_221_1_W0_addr),
    .W0_clk(mem_221_1_W0_clk),
    .W0_data(mem_221_1_W0_data),
    .W0_en(mem_221_1_W0_en),
    .W0_mask(mem_221_1_W0_mask)
  );
  split_mem_0_ext mem_221_2 (
    .R0_addr(mem_221_2_R0_addr),
    .R0_clk(mem_221_2_R0_clk),
    .R0_data(mem_221_2_R0_data),
    .R0_en(mem_221_2_R0_en),
    .W0_addr(mem_221_2_W0_addr),
    .W0_clk(mem_221_2_W0_clk),
    .W0_data(mem_221_2_W0_data),
    .W0_en(mem_221_2_W0_en),
    .W0_mask(mem_221_2_W0_mask)
  );
  split_mem_0_ext mem_221_3 (
    .R0_addr(mem_221_3_R0_addr),
    .R0_clk(mem_221_3_R0_clk),
    .R0_data(mem_221_3_R0_data),
    .R0_en(mem_221_3_R0_en),
    .W0_addr(mem_221_3_W0_addr),
    .W0_clk(mem_221_3_W0_clk),
    .W0_data(mem_221_3_W0_data),
    .W0_en(mem_221_3_W0_en),
    .W0_mask(mem_221_3_W0_mask)
  );
  split_mem_0_ext mem_221_4 (
    .R0_addr(mem_221_4_R0_addr),
    .R0_clk(mem_221_4_R0_clk),
    .R0_data(mem_221_4_R0_data),
    .R0_en(mem_221_4_R0_en),
    .W0_addr(mem_221_4_W0_addr),
    .W0_clk(mem_221_4_W0_clk),
    .W0_data(mem_221_4_W0_data),
    .W0_en(mem_221_4_W0_en),
    .W0_mask(mem_221_4_W0_mask)
  );
  split_mem_0_ext mem_221_5 (
    .R0_addr(mem_221_5_R0_addr),
    .R0_clk(mem_221_5_R0_clk),
    .R0_data(mem_221_5_R0_data),
    .R0_en(mem_221_5_R0_en),
    .W0_addr(mem_221_5_W0_addr),
    .W0_clk(mem_221_5_W0_clk),
    .W0_data(mem_221_5_W0_data),
    .W0_en(mem_221_5_W0_en),
    .W0_mask(mem_221_5_W0_mask)
  );
  split_mem_0_ext mem_221_6 (
    .R0_addr(mem_221_6_R0_addr),
    .R0_clk(mem_221_6_R0_clk),
    .R0_data(mem_221_6_R0_data),
    .R0_en(mem_221_6_R0_en),
    .W0_addr(mem_221_6_W0_addr),
    .W0_clk(mem_221_6_W0_clk),
    .W0_data(mem_221_6_W0_data),
    .W0_en(mem_221_6_W0_en),
    .W0_mask(mem_221_6_W0_mask)
  );
  split_mem_0_ext mem_221_7 (
    .R0_addr(mem_221_7_R0_addr),
    .R0_clk(mem_221_7_R0_clk),
    .R0_data(mem_221_7_R0_data),
    .R0_en(mem_221_7_R0_en),
    .W0_addr(mem_221_7_W0_addr),
    .W0_clk(mem_221_7_W0_clk),
    .W0_data(mem_221_7_W0_data),
    .W0_en(mem_221_7_W0_en),
    .W0_mask(mem_221_7_W0_mask)
  );
  split_mem_0_ext mem_222_0 (
    .R0_addr(mem_222_0_R0_addr),
    .R0_clk(mem_222_0_R0_clk),
    .R0_data(mem_222_0_R0_data),
    .R0_en(mem_222_0_R0_en),
    .W0_addr(mem_222_0_W0_addr),
    .W0_clk(mem_222_0_W0_clk),
    .W0_data(mem_222_0_W0_data),
    .W0_en(mem_222_0_W0_en),
    .W0_mask(mem_222_0_W0_mask)
  );
  split_mem_0_ext mem_222_1 (
    .R0_addr(mem_222_1_R0_addr),
    .R0_clk(mem_222_1_R0_clk),
    .R0_data(mem_222_1_R0_data),
    .R0_en(mem_222_1_R0_en),
    .W0_addr(mem_222_1_W0_addr),
    .W0_clk(mem_222_1_W0_clk),
    .W0_data(mem_222_1_W0_data),
    .W0_en(mem_222_1_W0_en),
    .W0_mask(mem_222_1_W0_mask)
  );
  split_mem_0_ext mem_222_2 (
    .R0_addr(mem_222_2_R0_addr),
    .R0_clk(mem_222_2_R0_clk),
    .R0_data(mem_222_2_R0_data),
    .R0_en(mem_222_2_R0_en),
    .W0_addr(mem_222_2_W0_addr),
    .W0_clk(mem_222_2_W0_clk),
    .W0_data(mem_222_2_W0_data),
    .W0_en(mem_222_2_W0_en),
    .W0_mask(mem_222_2_W0_mask)
  );
  split_mem_0_ext mem_222_3 (
    .R0_addr(mem_222_3_R0_addr),
    .R0_clk(mem_222_3_R0_clk),
    .R0_data(mem_222_3_R0_data),
    .R0_en(mem_222_3_R0_en),
    .W0_addr(mem_222_3_W0_addr),
    .W0_clk(mem_222_3_W0_clk),
    .W0_data(mem_222_3_W0_data),
    .W0_en(mem_222_3_W0_en),
    .W0_mask(mem_222_3_W0_mask)
  );
  split_mem_0_ext mem_222_4 (
    .R0_addr(mem_222_4_R0_addr),
    .R0_clk(mem_222_4_R0_clk),
    .R0_data(mem_222_4_R0_data),
    .R0_en(mem_222_4_R0_en),
    .W0_addr(mem_222_4_W0_addr),
    .W0_clk(mem_222_4_W0_clk),
    .W0_data(mem_222_4_W0_data),
    .W0_en(mem_222_4_W0_en),
    .W0_mask(mem_222_4_W0_mask)
  );
  split_mem_0_ext mem_222_5 (
    .R0_addr(mem_222_5_R0_addr),
    .R0_clk(mem_222_5_R0_clk),
    .R0_data(mem_222_5_R0_data),
    .R0_en(mem_222_5_R0_en),
    .W0_addr(mem_222_5_W0_addr),
    .W0_clk(mem_222_5_W0_clk),
    .W0_data(mem_222_5_W0_data),
    .W0_en(mem_222_5_W0_en),
    .W0_mask(mem_222_5_W0_mask)
  );
  split_mem_0_ext mem_222_6 (
    .R0_addr(mem_222_6_R0_addr),
    .R0_clk(mem_222_6_R0_clk),
    .R0_data(mem_222_6_R0_data),
    .R0_en(mem_222_6_R0_en),
    .W0_addr(mem_222_6_W0_addr),
    .W0_clk(mem_222_6_W0_clk),
    .W0_data(mem_222_6_W0_data),
    .W0_en(mem_222_6_W0_en),
    .W0_mask(mem_222_6_W0_mask)
  );
  split_mem_0_ext mem_222_7 (
    .R0_addr(mem_222_7_R0_addr),
    .R0_clk(mem_222_7_R0_clk),
    .R0_data(mem_222_7_R0_data),
    .R0_en(mem_222_7_R0_en),
    .W0_addr(mem_222_7_W0_addr),
    .W0_clk(mem_222_7_W0_clk),
    .W0_data(mem_222_7_W0_data),
    .W0_en(mem_222_7_W0_en),
    .W0_mask(mem_222_7_W0_mask)
  );
  split_mem_0_ext mem_223_0 (
    .R0_addr(mem_223_0_R0_addr),
    .R0_clk(mem_223_0_R0_clk),
    .R0_data(mem_223_0_R0_data),
    .R0_en(mem_223_0_R0_en),
    .W0_addr(mem_223_0_W0_addr),
    .W0_clk(mem_223_0_W0_clk),
    .W0_data(mem_223_0_W0_data),
    .W0_en(mem_223_0_W0_en),
    .W0_mask(mem_223_0_W0_mask)
  );
  split_mem_0_ext mem_223_1 (
    .R0_addr(mem_223_1_R0_addr),
    .R0_clk(mem_223_1_R0_clk),
    .R0_data(mem_223_1_R0_data),
    .R0_en(mem_223_1_R0_en),
    .W0_addr(mem_223_1_W0_addr),
    .W0_clk(mem_223_1_W0_clk),
    .W0_data(mem_223_1_W0_data),
    .W0_en(mem_223_1_W0_en),
    .W0_mask(mem_223_1_W0_mask)
  );
  split_mem_0_ext mem_223_2 (
    .R0_addr(mem_223_2_R0_addr),
    .R0_clk(mem_223_2_R0_clk),
    .R0_data(mem_223_2_R0_data),
    .R0_en(mem_223_2_R0_en),
    .W0_addr(mem_223_2_W0_addr),
    .W0_clk(mem_223_2_W0_clk),
    .W0_data(mem_223_2_W0_data),
    .W0_en(mem_223_2_W0_en),
    .W0_mask(mem_223_2_W0_mask)
  );
  split_mem_0_ext mem_223_3 (
    .R0_addr(mem_223_3_R0_addr),
    .R0_clk(mem_223_3_R0_clk),
    .R0_data(mem_223_3_R0_data),
    .R0_en(mem_223_3_R0_en),
    .W0_addr(mem_223_3_W0_addr),
    .W0_clk(mem_223_3_W0_clk),
    .W0_data(mem_223_3_W0_data),
    .W0_en(mem_223_3_W0_en),
    .W0_mask(mem_223_3_W0_mask)
  );
  split_mem_0_ext mem_223_4 (
    .R0_addr(mem_223_4_R0_addr),
    .R0_clk(mem_223_4_R0_clk),
    .R0_data(mem_223_4_R0_data),
    .R0_en(mem_223_4_R0_en),
    .W0_addr(mem_223_4_W0_addr),
    .W0_clk(mem_223_4_W0_clk),
    .W0_data(mem_223_4_W0_data),
    .W0_en(mem_223_4_W0_en),
    .W0_mask(mem_223_4_W0_mask)
  );
  split_mem_0_ext mem_223_5 (
    .R0_addr(mem_223_5_R0_addr),
    .R0_clk(mem_223_5_R0_clk),
    .R0_data(mem_223_5_R0_data),
    .R0_en(mem_223_5_R0_en),
    .W0_addr(mem_223_5_W0_addr),
    .W0_clk(mem_223_5_W0_clk),
    .W0_data(mem_223_5_W0_data),
    .W0_en(mem_223_5_W0_en),
    .W0_mask(mem_223_5_W0_mask)
  );
  split_mem_0_ext mem_223_6 (
    .R0_addr(mem_223_6_R0_addr),
    .R0_clk(mem_223_6_R0_clk),
    .R0_data(mem_223_6_R0_data),
    .R0_en(mem_223_6_R0_en),
    .W0_addr(mem_223_6_W0_addr),
    .W0_clk(mem_223_6_W0_clk),
    .W0_data(mem_223_6_W0_data),
    .W0_en(mem_223_6_W0_en),
    .W0_mask(mem_223_6_W0_mask)
  );
  split_mem_0_ext mem_223_7 (
    .R0_addr(mem_223_7_R0_addr),
    .R0_clk(mem_223_7_R0_clk),
    .R0_data(mem_223_7_R0_data),
    .R0_en(mem_223_7_R0_en),
    .W0_addr(mem_223_7_W0_addr),
    .W0_clk(mem_223_7_W0_clk),
    .W0_data(mem_223_7_W0_data),
    .W0_en(mem_223_7_W0_en),
    .W0_mask(mem_223_7_W0_mask)
  );
  split_mem_0_ext mem_224_0 (
    .R0_addr(mem_224_0_R0_addr),
    .R0_clk(mem_224_0_R0_clk),
    .R0_data(mem_224_0_R0_data),
    .R0_en(mem_224_0_R0_en),
    .W0_addr(mem_224_0_W0_addr),
    .W0_clk(mem_224_0_W0_clk),
    .W0_data(mem_224_0_W0_data),
    .W0_en(mem_224_0_W0_en),
    .W0_mask(mem_224_0_W0_mask)
  );
  split_mem_0_ext mem_224_1 (
    .R0_addr(mem_224_1_R0_addr),
    .R0_clk(mem_224_1_R0_clk),
    .R0_data(mem_224_1_R0_data),
    .R0_en(mem_224_1_R0_en),
    .W0_addr(mem_224_1_W0_addr),
    .W0_clk(mem_224_1_W0_clk),
    .W0_data(mem_224_1_W0_data),
    .W0_en(mem_224_1_W0_en),
    .W0_mask(mem_224_1_W0_mask)
  );
  split_mem_0_ext mem_224_2 (
    .R0_addr(mem_224_2_R0_addr),
    .R0_clk(mem_224_2_R0_clk),
    .R0_data(mem_224_2_R0_data),
    .R0_en(mem_224_2_R0_en),
    .W0_addr(mem_224_2_W0_addr),
    .W0_clk(mem_224_2_W0_clk),
    .W0_data(mem_224_2_W0_data),
    .W0_en(mem_224_2_W0_en),
    .W0_mask(mem_224_2_W0_mask)
  );
  split_mem_0_ext mem_224_3 (
    .R0_addr(mem_224_3_R0_addr),
    .R0_clk(mem_224_3_R0_clk),
    .R0_data(mem_224_3_R0_data),
    .R0_en(mem_224_3_R0_en),
    .W0_addr(mem_224_3_W0_addr),
    .W0_clk(mem_224_3_W0_clk),
    .W0_data(mem_224_3_W0_data),
    .W0_en(mem_224_3_W0_en),
    .W0_mask(mem_224_3_W0_mask)
  );
  split_mem_0_ext mem_224_4 (
    .R0_addr(mem_224_4_R0_addr),
    .R0_clk(mem_224_4_R0_clk),
    .R0_data(mem_224_4_R0_data),
    .R0_en(mem_224_4_R0_en),
    .W0_addr(mem_224_4_W0_addr),
    .W0_clk(mem_224_4_W0_clk),
    .W0_data(mem_224_4_W0_data),
    .W0_en(mem_224_4_W0_en),
    .W0_mask(mem_224_4_W0_mask)
  );
  split_mem_0_ext mem_224_5 (
    .R0_addr(mem_224_5_R0_addr),
    .R0_clk(mem_224_5_R0_clk),
    .R0_data(mem_224_5_R0_data),
    .R0_en(mem_224_5_R0_en),
    .W0_addr(mem_224_5_W0_addr),
    .W0_clk(mem_224_5_W0_clk),
    .W0_data(mem_224_5_W0_data),
    .W0_en(mem_224_5_W0_en),
    .W0_mask(mem_224_5_W0_mask)
  );
  split_mem_0_ext mem_224_6 (
    .R0_addr(mem_224_6_R0_addr),
    .R0_clk(mem_224_6_R0_clk),
    .R0_data(mem_224_6_R0_data),
    .R0_en(mem_224_6_R0_en),
    .W0_addr(mem_224_6_W0_addr),
    .W0_clk(mem_224_6_W0_clk),
    .W0_data(mem_224_6_W0_data),
    .W0_en(mem_224_6_W0_en),
    .W0_mask(mem_224_6_W0_mask)
  );
  split_mem_0_ext mem_224_7 (
    .R0_addr(mem_224_7_R0_addr),
    .R0_clk(mem_224_7_R0_clk),
    .R0_data(mem_224_7_R0_data),
    .R0_en(mem_224_7_R0_en),
    .W0_addr(mem_224_7_W0_addr),
    .W0_clk(mem_224_7_W0_clk),
    .W0_data(mem_224_7_W0_data),
    .W0_en(mem_224_7_W0_en),
    .W0_mask(mem_224_7_W0_mask)
  );
  split_mem_0_ext mem_225_0 (
    .R0_addr(mem_225_0_R0_addr),
    .R0_clk(mem_225_0_R0_clk),
    .R0_data(mem_225_0_R0_data),
    .R0_en(mem_225_0_R0_en),
    .W0_addr(mem_225_0_W0_addr),
    .W0_clk(mem_225_0_W0_clk),
    .W0_data(mem_225_0_W0_data),
    .W0_en(mem_225_0_W0_en),
    .W0_mask(mem_225_0_W0_mask)
  );
  split_mem_0_ext mem_225_1 (
    .R0_addr(mem_225_1_R0_addr),
    .R0_clk(mem_225_1_R0_clk),
    .R0_data(mem_225_1_R0_data),
    .R0_en(mem_225_1_R0_en),
    .W0_addr(mem_225_1_W0_addr),
    .W0_clk(mem_225_1_W0_clk),
    .W0_data(mem_225_1_W0_data),
    .W0_en(mem_225_1_W0_en),
    .W0_mask(mem_225_1_W0_mask)
  );
  split_mem_0_ext mem_225_2 (
    .R0_addr(mem_225_2_R0_addr),
    .R0_clk(mem_225_2_R0_clk),
    .R0_data(mem_225_2_R0_data),
    .R0_en(mem_225_2_R0_en),
    .W0_addr(mem_225_2_W0_addr),
    .W0_clk(mem_225_2_W0_clk),
    .W0_data(mem_225_2_W0_data),
    .W0_en(mem_225_2_W0_en),
    .W0_mask(mem_225_2_W0_mask)
  );
  split_mem_0_ext mem_225_3 (
    .R0_addr(mem_225_3_R0_addr),
    .R0_clk(mem_225_3_R0_clk),
    .R0_data(mem_225_3_R0_data),
    .R0_en(mem_225_3_R0_en),
    .W0_addr(mem_225_3_W0_addr),
    .W0_clk(mem_225_3_W0_clk),
    .W0_data(mem_225_3_W0_data),
    .W0_en(mem_225_3_W0_en),
    .W0_mask(mem_225_3_W0_mask)
  );
  split_mem_0_ext mem_225_4 (
    .R0_addr(mem_225_4_R0_addr),
    .R0_clk(mem_225_4_R0_clk),
    .R0_data(mem_225_4_R0_data),
    .R0_en(mem_225_4_R0_en),
    .W0_addr(mem_225_4_W0_addr),
    .W0_clk(mem_225_4_W0_clk),
    .W0_data(mem_225_4_W0_data),
    .W0_en(mem_225_4_W0_en),
    .W0_mask(mem_225_4_W0_mask)
  );
  split_mem_0_ext mem_225_5 (
    .R0_addr(mem_225_5_R0_addr),
    .R0_clk(mem_225_5_R0_clk),
    .R0_data(mem_225_5_R0_data),
    .R0_en(mem_225_5_R0_en),
    .W0_addr(mem_225_5_W0_addr),
    .W0_clk(mem_225_5_W0_clk),
    .W0_data(mem_225_5_W0_data),
    .W0_en(mem_225_5_W0_en),
    .W0_mask(mem_225_5_W0_mask)
  );
  split_mem_0_ext mem_225_6 (
    .R0_addr(mem_225_6_R0_addr),
    .R0_clk(mem_225_6_R0_clk),
    .R0_data(mem_225_6_R0_data),
    .R0_en(mem_225_6_R0_en),
    .W0_addr(mem_225_6_W0_addr),
    .W0_clk(mem_225_6_W0_clk),
    .W0_data(mem_225_6_W0_data),
    .W0_en(mem_225_6_W0_en),
    .W0_mask(mem_225_6_W0_mask)
  );
  split_mem_0_ext mem_225_7 (
    .R0_addr(mem_225_7_R0_addr),
    .R0_clk(mem_225_7_R0_clk),
    .R0_data(mem_225_7_R0_data),
    .R0_en(mem_225_7_R0_en),
    .W0_addr(mem_225_7_W0_addr),
    .W0_clk(mem_225_7_W0_clk),
    .W0_data(mem_225_7_W0_data),
    .W0_en(mem_225_7_W0_en),
    .W0_mask(mem_225_7_W0_mask)
  );
  split_mem_0_ext mem_226_0 (
    .R0_addr(mem_226_0_R0_addr),
    .R0_clk(mem_226_0_R0_clk),
    .R0_data(mem_226_0_R0_data),
    .R0_en(mem_226_0_R0_en),
    .W0_addr(mem_226_0_W0_addr),
    .W0_clk(mem_226_0_W0_clk),
    .W0_data(mem_226_0_W0_data),
    .W0_en(mem_226_0_W0_en),
    .W0_mask(mem_226_0_W0_mask)
  );
  split_mem_0_ext mem_226_1 (
    .R0_addr(mem_226_1_R0_addr),
    .R0_clk(mem_226_1_R0_clk),
    .R0_data(mem_226_1_R0_data),
    .R0_en(mem_226_1_R0_en),
    .W0_addr(mem_226_1_W0_addr),
    .W0_clk(mem_226_1_W0_clk),
    .W0_data(mem_226_1_W0_data),
    .W0_en(mem_226_1_W0_en),
    .W0_mask(mem_226_1_W0_mask)
  );
  split_mem_0_ext mem_226_2 (
    .R0_addr(mem_226_2_R0_addr),
    .R0_clk(mem_226_2_R0_clk),
    .R0_data(mem_226_2_R0_data),
    .R0_en(mem_226_2_R0_en),
    .W0_addr(mem_226_2_W0_addr),
    .W0_clk(mem_226_2_W0_clk),
    .W0_data(mem_226_2_W0_data),
    .W0_en(mem_226_2_W0_en),
    .W0_mask(mem_226_2_W0_mask)
  );
  split_mem_0_ext mem_226_3 (
    .R0_addr(mem_226_3_R0_addr),
    .R0_clk(mem_226_3_R0_clk),
    .R0_data(mem_226_3_R0_data),
    .R0_en(mem_226_3_R0_en),
    .W0_addr(mem_226_3_W0_addr),
    .W0_clk(mem_226_3_W0_clk),
    .W0_data(mem_226_3_W0_data),
    .W0_en(mem_226_3_W0_en),
    .W0_mask(mem_226_3_W0_mask)
  );
  split_mem_0_ext mem_226_4 (
    .R0_addr(mem_226_4_R0_addr),
    .R0_clk(mem_226_4_R0_clk),
    .R0_data(mem_226_4_R0_data),
    .R0_en(mem_226_4_R0_en),
    .W0_addr(mem_226_4_W0_addr),
    .W0_clk(mem_226_4_W0_clk),
    .W0_data(mem_226_4_W0_data),
    .W0_en(mem_226_4_W0_en),
    .W0_mask(mem_226_4_W0_mask)
  );
  split_mem_0_ext mem_226_5 (
    .R0_addr(mem_226_5_R0_addr),
    .R0_clk(mem_226_5_R0_clk),
    .R0_data(mem_226_5_R0_data),
    .R0_en(mem_226_5_R0_en),
    .W0_addr(mem_226_5_W0_addr),
    .W0_clk(mem_226_5_W0_clk),
    .W0_data(mem_226_5_W0_data),
    .W0_en(mem_226_5_W0_en),
    .W0_mask(mem_226_5_W0_mask)
  );
  split_mem_0_ext mem_226_6 (
    .R0_addr(mem_226_6_R0_addr),
    .R0_clk(mem_226_6_R0_clk),
    .R0_data(mem_226_6_R0_data),
    .R0_en(mem_226_6_R0_en),
    .W0_addr(mem_226_6_W0_addr),
    .W0_clk(mem_226_6_W0_clk),
    .W0_data(mem_226_6_W0_data),
    .W0_en(mem_226_6_W0_en),
    .W0_mask(mem_226_6_W0_mask)
  );
  split_mem_0_ext mem_226_7 (
    .R0_addr(mem_226_7_R0_addr),
    .R0_clk(mem_226_7_R0_clk),
    .R0_data(mem_226_7_R0_data),
    .R0_en(mem_226_7_R0_en),
    .W0_addr(mem_226_7_W0_addr),
    .W0_clk(mem_226_7_W0_clk),
    .W0_data(mem_226_7_W0_data),
    .W0_en(mem_226_7_W0_en),
    .W0_mask(mem_226_7_W0_mask)
  );
  split_mem_0_ext mem_227_0 (
    .R0_addr(mem_227_0_R0_addr),
    .R0_clk(mem_227_0_R0_clk),
    .R0_data(mem_227_0_R0_data),
    .R0_en(mem_227_0_R0_en),
    .W0_addr(mem_227_0_W0_addr),
    .W0_clk(mem_227_0_W0_clk),
    .W0_data(mem_227_0_W0_data),
    .W0_en(mem_227_0_W0_en),
    .W0_mask(mem_227_0_W0_mask)
  );
  split_mem_0_ext mem_227_1 (
    .R0_addr(mem_227_1_R0_addr),
    .R0_clk(mem_227_1_R0_clk),
    .R0_data(mem_227_1_R0_data),
    .R0_en(mem_227_1_R0_en),
    .W0_addr(mem_227_1_W0_addr),
    .W0_clk(mem_227_1_W0_clk),
    .W0_data(mem_227_1_W0_data),
    .W0_en(mem_227_1_W0_en),
    .W0_mask(mem_227_1_W0_mask)
  );
  split_mem_0_ext mem_227_2 (
    .R0_addr(mem_227_2_R0_addr),
    .R0_clk(mem_227_2_R0_clk),
    .R0_data(mem_227_2_R0_data),
    .R0_en(mem_227_2_R0_en),
    .W0_addr(mem_227_2_W0_addr),
    .W0_clk(mem_227_2_W0_clk),
    .W0_data(mem_227_2_W0_data),
    .W0_en(mem_227_2_W0_en),
    .W0_mask(mem_227_2_W0_mask)
  );
  split_mem_0_ext mem_227_3 (
    .R0_addr(mem_227_3_R0_addr),
    .R0_clk(mem_227_3_R0_clk),
    .R0_data(mem_227_3_R0_data),
    .R0_en(mem_227_3_R0_en),
    .W0_addr(mem_227_3_W0_addr),
    .W0_clk(mem_227_3_W0_clk),
    .W0_data(mem_227_3_W0_data),
    .W0_en(mem_227_3_W0_en),
    .W0_mask(mem_227_3_W0_mask)
  );
  split_mem_0_ext mem_227_4 (
    .R0_addr(mem_227_4_R0_addr),
    .R0_clk(mem_227_4_R0_clk),
    .R0_data(mem_227_4_R0_data),
    .R0_en(mem_227_4_R0_en),
    .W0_addr(mem_227_4_W0_addr),
    .W0_clk(mem_227_4_W0_clk),
    .W0_data(mem_227_4_W0_data),
    .W0_en(mem_227_4_W0_en),
    .W0_mask(mem_227_4_W0_mask)
  );
  split_mem_0_ext mem_227_5 (
    .R0_addr(mem_227_5_R0_addr),
    .R0_clk(mem_227_5_R0_clk),
    .R0_data(mem_227_5_R0_data),
    .R0_en(mem_227_5_R0_en),
    .W0_addr(mem_227_5_W0_addr),
    .W0_clk(mem_227_5_W0_clk),
    .W0_data(mem_227_5_W0_data),
    .W0_en(mem_227_5_W0_en),
    .W0_mask(mem_227_5_W0_mask)
  );
  split_mem_0_ext mem_227_6 (
    .R0_addr(mem_227_6_R0_addr),
    .R0_clk(mem_227_6_R0_clk),
    .R0_data(mem_227_6_R0_data),
    .R0_en(mem_227_6_R0_en),
    .W0_addr(mem_227_6_W0_addr),
    .W0_clk(mem_227_6_W0_clk),
    .W0_data(mem_227_6_W0_data),
    .W0_en(mem_227_6_W0_en),
    .W0_mask(mem_227_6_W0_mask)
  );
  split_mem_0_ext mem_227_7 (
    .R0_addr(mem_227_7_R0_addr),
    .R0_clk(mem_227_7_R0_clk),
    .R0_data(mem_227_7_R0_data),
    .R0_en(mem_227_7_R0_en),
    .W0_addr(mem_227_7_W0_addr),
    .W0_clk(mem_227_7_W0_clk),
    .W0_data(mem_227_7_W0_data),
    .W0_en(mem_227_7_W0_en),
    .W0_mask(mem_227_7_W0_mask)
  );
  split_mem_0_ext mem_228_0 (
    .R0_addr(mem_228_0_R0_addr),
    .R0_clk(mem_228_0_R0_clk),
    .R0_data(mem_228_0_R0_data),
    .R0_en(mem_228_0_R0_en),
    .W0_addr(mem_228_0_W0_addr),
    .W0_clk(mem_228_0_W0_clk),
    .W0_data(mem_228_0_W0_data),
    .W0_en(mem_228_0_W0_en),
    .W0_mask(mem_228_0_W0_mask)
  );
  split_mem_0_ext mem_228_1 (
    .R0_addr(mem_228_1_R0_addr),
    .R0_clk(mem_228_1_R0_clk),
    .R0_data(mem_228_1_R0_data),
    .R0_en(mem_228_1_R0_en),
    .W0_addr(mem_228_1_W0_addr),
    .W0_clk(mem_228_1_W0_clk),
    .W0_data(mem_228_1_W0_data),
    .W0_en(mem_228_1_W0_en),
    .W0_mask(mem_228_1_W0_mask)
  );
  split_mem_0_ext mem_228_2 (
    .R0_addr(mem_228_2_R0_addr),
    .R0_clk(mem_228_2_R0_clk),
    .R0_data(mem_228_2_R0_data),
    .R0_en(mem_228_2_R0_en),
    .W0_addr(mem_228_2_W0_addr),
    .W0_clk(mem_228_2_W0_clk),
    .W0_data(mem_228_2_W0_data),
    .W0_en(mem_228_2_W0_en),
    .W0_mask(mem_228_2_W0_mask)
  );
  split_mem_0_ext mem_228_3 (
    .R0_addr(mem_228_3_R0_addr),
    .R0_clk(mem_228_3_R0_clk),
    .R0_data(mem_228_3_R0_data),
    .R0_en(mem_228_3_R0_en),
    .W0_addr(mem_228_3_W0_addr),
    .W0_clk(mem_228_3_W0_clk),
    .W0_data(mem_228_3_W0_data),
    .W0_en(mem_228_3_W0_en),
    .W0_mask(mem_228_3_W0_mask)
  );
  split_mem_0_ext mem_228_4 (
    .R0_addr(mem_228_4_R0_addr),
    .R0_clk(mem_228_4_R0_clk),
    .R0_data(mem_228_4_R0_data),
    .R0_en(mem_228_4_R0_en),
    .W0_addr(mem_228_4_W0_addr),
    .W0_clk(mem_228_4_W0_clk),
    .W0_data(mem_228_4_W0_data),
    .W0_en(mem_228_4_W0_en),
    .W0_mask(mem_228_4_W0_mask)
  );
  split_mem_0_ext mem_228_5 (
    .R0_addr(mem_228_5_R0_addr),
    .R0_clk(mem_228_5_R0_clk),
    .R0_data(mem_228_5_R0_data),
    .R0_en(mem_228_5_R0_en),
    .W0_addr(mem_228_5_W0_addr),
    .W0_clk(mem_228_5_W0_clk),
    .W0_data(mem_228_5_W0_data),
    .W0_en(mem_228_5_W0_en),
    .W0_mask(mem_228_5_W0_mask)
  );
  split_mem_0_ext mem_228_6 (
    .R0_addr(mem_228_6_R0_addr),
    .R0_clk(mem_228_6_R0_clk),
    .R0_data(mem_228_6_R0_data),
    .R0_en(mem_228_6_R0_en),
    .W0_addr(mem_228_6_W0_addr),
    .W0_clk(mem_228_6_W0_clk),
    .W0_data(mem_228_6_W0_data),
    .W0_en(mem_228_6_W0_en),
    .W0_mask(mem_228_6_W0_mask)
  );
  split_mem_0_ext mem_228_7 (
    .R0_addr(mem_228_7_R0_addr),
    .R0_clk(mem_228_7_R0_clk),
    .R0_data(mem_228_7_R0_data),
    .R0_en(mem_228_7_R0_en),
    .W0_addr(mem_228_7_W0_addr),
    .W0_clk(mem_228_7_W0_clk),
    .W0_data(mem_228_7_W0_data),
    .W0_en(mem_228_7_W0_en),
    .W0_mask(mem_228_7_W0_mask)
  );
  split_mem_0_ext mem_229_0 (
    .R0_addr(mem_229_0_R0_addr),
    .R0_clk(mem_229_0_R0_clk),
    .R0_data(mem_229_0_R0_data),
    .R0_en(mem_229_0_R0_en),
    .W0_addr(mem_229_0_W0_addr),
    .W0_clk(mem_229_0_W0_clk),
    .W0_data(mem_229_0_W0_data),
    .W0_en(mem_229_0_W0_en),
    .W0_mask(mem_229_0_W0_mask)
  );
  split_mem_0_ext mem_229_1 (
    .R0_addr(mem_229_1_R0_addr),
    .R0_clk(mem_229_1_R0_clk),
    .R0_data(mem_229_1_R0_data),
    .R0_en(mem_229_1_R0_en),
    .W0_addr(mem_229_1_W0_addr),
    .W0_clk(mem_229_1_W0_clk),
    .W0_data(mem_229_1_W0_data),
    .W0_en(mem_229_1_W0_en),
    .W0_mask(mem_229_1_W0_mask)
  );
  split_mem_0_ext mem_229_2 (
    .R0_addr(mem_229_2_R0_addr),
    .R0_clk(mem_229_2_R0_clk),
    .R0_data(mem_229_2_R0_data),
    .R0_en(mem_229_2_R0_en),
    .W0_addr(mem_229_2_W0_addr),
    .W0_clk(mem_229_2_W0_clk),
    .W0_data(mem_229_2_W0_data),
    .W0_en(mem_229_2_W0_en),
    .W0_mask(mem_229_2_W0_mask)
  );
  split_mem_0_ext mem_229_3 (
    .R0_addr(mem_229_3_R0_addr),
    .R0_clk(mem_229_3_R0_clk),
    .R0_data(mem_229_3_R0_data),
    .R0_en(mem_229_3_R0_en),
    .W0_addr(mem_229_3_W0_addr),
    .W0_clk(mem_229_3_W0_clk),
    .W0_data(mem_229_3_W0_data),
    .W0_en(mem_229_3_W0_en),
    .W0_mask(mem_229_3_W0_mask)
  );
  split_mem_0_ext mem_229_4 (
    .R0_addr(mem_229_4_R0_addr),
    .R0_clk(mem_229_4_R0_clk),
    .R0_data(mem_229_4_R0_data),
    .R0_en(mem_229_4_R0_en),
    .W0_addr(mem_229_4_W0_addr),
    .W0_clk(mem_229_4_W0_clk),
    .W0_data(mem_229_4_W0_data),
    .W0_en(mem_229_4_W0_en),
    .W0_mask(mem_229_4_W0_mask)
  );
  split_mem_0_ext mem_229_5 (
    .R0_addr(mem_229_5_R0_addr),
    .R0_clk(mem_229_5_R0_clk),
    .R0_data(mem_229_5_R0_data),
    .R0_en(mem_229_5_R0_en),
    .W0_addr(mem_229_5_W0_addr),
    .W0_clk(mem_229_5_W0_clk),
    .W0_data(mem_229_5_W0_data),
    .W0_en(mem_229_5_W0_en),
    .W0_mask(mem_229_5_W0_mask)
  );
  split_mem_0_ext mem_229_6 (
    .R0_addr(mem_229_6_R0_addr),
    .R0_clk(mem_229_6_R0_clk),
    .R0_data(mem_229_6_R0_data),
    .R0_en(mem_229_6_R0_en),
    .W0_addr(mem_229_6_W0_addr),
    .W0_clk(mem_229_6_W0_clk),
    .W0_data(mem_229_6_W0_data),
    .W0_en(mem_229_6_W0_en),
    .W0_mask(mem_229_6_W0_mask)
  );
  split_mem_0_ext mem_229_7 (
    .R0_addr(mem_229_7_R0_addr),
    .R0_clk(mem_229_7_R0_clk),
    .R0_data(mem_229_7_R0_data),
    .R0_en(mem_229_7_R0_en),
    .W0_addr(mem_229_7_W0_addr),
    .W0_clk(mem_229_7_W0_clk),
    .W0_data(mem_229_7_W0_data),
    .W0_en(mem_229_7_W0_en),
    .W0_mask(mem_229_7_W0_mask)
  );
  split_mem_0_ext mem_230_0 (
    .R0_addr(mem_230_0_R0_addr),
    .R0_clk(mem_230_0_R0_clk),
    .R0_data(mem_230_0_R0_data),
    .R0_en(mem_230_0_R0_en),
    .W0_addr(mem_230_0_W0_addr),
    .W0_clk(mem_230_0_W0_clk),
    .W0_data(mem_230_0_W0_data),
    .W0_en(mem_230_0_W0_en),
    .W0_mask(mem_230_0_W0_mask)
  );
  split_mem_0_ext mem_230_1 (
    .R0_addr(mem_230_1_R0_addr),
    .R0_clk(mem_230_1_R0_clk),
    .R0_data(mem_230_1_R0_data),
    .R0_en(mem_230_1_R0_en),
    .W0_addr(mem_230_1_W0_addr),
    .W0_clk(mem_230_1_W0_clk),
    .W0_data(mem_230_1_W0_data),
    .W0_en(mem_230_1_W0_en),
    .W0_mask(mem_230_1_W0_mask)
  );
  split_mem_0_ext mem_230_2 (
    .R0_addr(mem_230_2_R0_addr),
    .R0_clk(mem_230_2_R0_clk),
    .R0_data(mem_230_2_R0_data),
    .R0_en(mem_230_2_R0_en),
    .W0_addr(mem_230_2_W0_addr),
    .W0_clk(mem_230_2_W0_clk),
    .W0_data(mem_230_2_W0_data),
    .W0_en(mem_230_2_W0_en),
    .W0_mask(mem_230_2_W0_mask)
  );
  split_mem_0_ext mem_230_3 (
    .R0_addr(mem_230_3_R0_addr),
    .R0_clk(mem_230_3_R0_clk),
    .R0_data(mem_230_3_R0_data),
    .R0_en(mem_230_3_R0_en),
    .W0_addr(mem_230_3_W0_addr),
    .W0_clk(mem_230_3_W0_clk),
    .W0_data(mem_230_3_W0_data),
    .W0_en(mem_230_3_W0_en),
    .W0_mask(mem_230_3_W0_mask)
  );
  split_mem_0_ext mem_230_4 (
    .R0_addr(mem_230_4_R0_addr),
    .R0_clk(mem_230_4_R0_clk),
    .R0_data(mem_230_4_R0_data),
    .R0_en(mem_230_4_R0_en),
    .W0_addr(mem_230_4_W0_addr),
    .W0_clk(mem_230_4_W0_clk),
    .W0_data(mem_230_4_W0_data),
    .W0_en(mem_230_4_W0_en),
    .W0_mask(mem_230_4_W0_mask)
  );
  split_mem_0_ext mem_230_5 (
    .R0_addr(mem_230_5_R0_addr),
    .R0_clk(mem_230_5_R0_clk),
    .R0_data(mem_230_5_R0_data),
    .R0_en(mem_230_5_R0_en),
    .W0_addr(mem_230_5_W0_addr),
    .W0_clk(mem_230_5_W0_clk),
    .W0_data(mem_230_5_W0_data),
    .W0_en(mem_230_5_W0_en),
    .W0_mask(mem_230_5_W0_mask)
  );
  split_mem_0_ext mem_230_6 (
    .R0_addr(mem_230_6_R0_addr),
    .R0_clk(mem_230_6_R0_clk),
    .R0_data(mem_230_6_R0_data),
    .R0_en(mem_230_6_R0_en),
    .W0_addr(mem_230_6_W0_addr),
    .W0_clk(mem_230_6_W0_clk),
    .W0_data(mem_230_6_W0_data),
    .W0_en(mem_230_6_W0_en),
    .W0_mask(mem_230_6_W0_mask)
  );
  split_mem_0_ext mem_230_7 (
    .R0_addr(mem_230_7_R0_addr),
    .R0_clk(mem_230_7_R0_clk),
    .R0_data(mem_230_7_R0_data),
    .R0_en(mem_230_7_R0_en),
    .W0_addr(mem_230_7_W0_addr),
    .W0_clk(mem_230_7_W0_clk),
    .W0_data(mem_230_7_W0_data),
    .W0_en(mem_230_7_W0_en),
    .W0_mask(mem_230_7_W0_mask)
  );
  split_mem_0_ext mem_231_0 (
    .R0_addr(mem_231_0_R0_addr),
    .R0_clk(mem_231_0_R0_clk),
    .R0_data(mem_231_0_R0_data),
    .R0_en(mem_231_0_R0_en),
    .W0_addr(mem_231_0_W0_addr),
    .W0_clk(mem_231_0_W0_clk),
    .W0_data(mem_231_0_W0_data),
    .W0_en(mem_231_0_W0_en),
    .W0_mask(mem_231_0_W0_mask)
  );
  split_mem_0_ext mem_231_1 (
    .R0_addr(mem_231_1_R0_addr),
    .R0_clk(mem_231_1_R0_clk),
    .R0_data(mem_231_1_R0_data),
    .R0_en(mem_231_1_R0_en),
    .W0_addr(mem_231_1_W0_addr),
    .W0_clk(mem_231_1_W0_clk),
    .W0_data(mem_231_1_W0_data),
    .W0_en(mem_231_1_W0_en),
    .W0_mask(mem_231_1_W0_mask)
  );
  split_mem_0_ext mem_231_2 (
    .R0_addr(mem_231_2_R0_addr),
    .R0_clk(mem_231_2_R0_clk),
    .R0_data(mem_231_2_R0_data),
    .R0_en(mem_231_2_R0_en),
    .W0_addr(mem_231_2_W0_addr),
    .W0_clk(mem_231_2_W0_clk),
    .W0_data(mem_231_2_W0_data),
    .W0_en(mem_231_2_W0_en),
    .W0_mask(mem_231_2_W0_mask)
  );
  split_mem_0_ext mem_231_3 (
    .R0_addr(mem_231_3_R0_addr),
    .R0_clk(mem_231_3_R0_clk),
    .R0_data(mem_231_3_R0_data),
    .R0_en(mem_231_3_R0_en),
    .W0_addr(mem_231_3_W0_addr),
    .W0_clk(mem_231_3_W0_clk),
    .W0_data(mem_231_3_W0_data),
    .W0_en(mem_231_3_W0_en),
    .W0_mask(mem_231_3_W0_mask)
  );
  split_mem_0_ext mem_231_4 (
    .R0_addr(mem_231_4_R0_addr),
    .R0_clk(mem_231_4_R0_clk),
    .R0_data(mem_231_4_R0_data),
    .R0_en(mem_231_4_R0_en),
    .W0_addr(mem_231_4_W0_addr),
    .W0_clk(mem_231_4_W0_clk),
    .W0_data(mem_231_4_W0_data),
    .W0_en(mem_231_4_W0_en),
    .W0_mask(mem_231_4_W0_mask)
  );
  split_mem_0_ext mem_231_5 (
    .R0_addr(mem_231_5_R0_addr),
    .R0_clk(mem_231_5_R0_clk),
    .R0_data(mem_231_5_R0_data),
    .R0_en(mem_231_5_R0_en),
    .W0_addr(mem_231_5_W0_addr),
    .W0_clk(mem_231_5_W0_clk),
    .W0_data(mem_231_5_W0_data),
    .W0_en(mem_231_5_W0_en),
    .W0_mask(mem_231_5_W0_mask)
  );
  split_mem_0_ext mem_231_6 (
    .R0_addr(mem_231_6_R0_addr),
    .R0_clk(mem_231_6_R0_clk),
    .R0_data(mem_231_6_R0_data),
    .R0_en(mem_231_6_R0_en),
    .W0_addr(mem_231_6_W0_addr),
    .W0_clk(mem_231_6_W0_clk),
    .W0_data(mem_231_6_W0_data),
    .W0_en(mem_231_6_W0_en),
    .W0_mask(mem_231_6_W0_mask)
  );
  split_mem_0_ext mem_231_7 (
    .R0_addr(mem_231_7_R0_addr),
    .R0_clk(mem_231_7_R0_clk),
    .R0_data(mem_231_7_R0_data),
    .R0_en(mem_231_7_R0_en),
    .W0_addr(mem_231_7_W0_addr),
    .W0_clk(mem_231_7_W0_clk),
    .W0_data(mem_231_7_W0_data),
    .W0_en(mem_231_7_W0_en),
    .W0_mask(mem_231_7_W0_mask)
  );
  split_mem_0_ext mem_232_0 (
    .R0_addr(mem_232_0_R0_addr),
    .R0_clk(mem_232_0_R0_clk),
    .R0_data(mem_232_0_R0_data),
    .R0_en(mem_232_0_R0_en),
    .W0_addr(mem_232_0_W0_addr),
    .W0_clk(mem_232_0_W0_clk),
    .W0_data(mem_232_0_W0_data),
    .W0_en(mem_232_0_W0_en),
    .W0_mask(mem_232_0_W0_mask)
  );
  split_mem_0_ext mem_232_1 (
    .R0_addr(mem_232_1_R0_addr),
    .R0_clk(mem_232_1_R0_clk),
    .R0_data(mem_232_1_R0_data),
    .R0_en(mem_232_1_R0_en),
    .W0_addr(mem_232_1_W0_addr),
    .W0_clk(mem_232_1_W0_clk),
    .W0_data(mem_232_1_W0_data),
    .W0_en(mem_232_1_W0_en),
    .W0_mask(mem_232_1_W0_mask)
  );
  split_mem_0_ext mem_232_2 (
    .R0_addr(mem_232_2_R0_addr),
    .R0_clk(mem_232_2_R0_clk),
    .R0_data(mem_232_2_R0_data),
    .R0_en(mem_232_2_R0_en),
    .W0_addr(mem_232_2_W0_addr),
    .W0_clk(mem_232_2_W0_clk),
    .W0_data(mem_232_2_W0_data),
    .W0_en(mem_232_2_W0_en),
    .W0_mask(mem_232_2_W0_mask)
  );
  split_mem_0_ext mem_232_3 (
    .R0_addr(mem_232_3_R0_addr),
    .R0_clk(mem_232_3_R0_clk),
    .R0_data(mem_232_3_R0_data),
    .R0_en(mem_232_3_R0_en),
    .W0_addr(mem_232_3_W0_addr),
    .W0_clk(mem_232_3_W0_clk),
    .W0_data(mem_232_3_W0_data),
    .W0_en(mem_232_3_W0_en),
    .W0_mask(mem_232_3_W0_mask)
  );
  split_mem_0_ext mem_232_4 (
    .R0_addr(mem_232_4_R0_addr),
    .R0_clk(mem_232_4_R0_clk),
    .R0_data(mem_232_4_R0_data),
    .R0_en(mem_232_4_R0_en),
    .W0_addr(mem_232_4_W0_addr),
    .W0_clk(mem_232_4_W0_clk),
    .W0_data(mem_232_4_W0_data),
    .W0_en(mem_232_4_W0_en),
    .W0_mask(mem_232_4_W0_mask)
  );
  split_mem_0_ext mem_232_5 (
    .R0_addr(mem_232_5_R0_addr),
    .R0_clk(mem_232_5_R0_clk),
    .R0_data(mem_232_5_R0_data),
    .R0_en(mem_232_5_R0_en),
    .W0_addr(mem_232_5_W0_addr),
    .W0_clk(mem_232_5_W0_clk),
    .W0_data(mem_232_5_W0_data),
    .W0_en(mem_232_5_W0_en),
    .W0_mask(mem_232_5_W0_mask)
  );
  split_mem_0_ext mem_232_6 (
    .R0_addr(mem_232_6_R0_addr),
    .R0_clk(mem_232_6_R0_clk),
    .R0_data(mem_232_6_R0_data),
    .R0_en(mem_232_6_R0_en),
    .W0_addr(mem_232_6_W0_addr),
    .W0_clk(mem_232_6_W0_clk),
    .W0_data(mem_232_6_W0_data),
    .W0_en(mem_232_6_W0_en),
    .W0_mask(mem_232_6_W0_mask)
  );
  split_mem_0_ext mem_232_7 (
    .R0_addr(mem_232_7_R0_addr),
    .R0_clk(mem_232_7_R0_clk),
    .R0_data(mem_232_7_R0_data),
    .R0_en(mem_232_7_R0_en),
    .W0_addr(mem_232_7_W0_addr),
    .W0_clk(mem_232_7_W0_clk),
    .W0_data(mem_232_7_W0_data),
    .W0_en(mem_232_7_W0_en),
    .W0_mask(mem_232_7_W0_mask)
  );
  split_mem_0_ext mem_233_0 (
    .R0_addr(mem_233_0_R0_addr),
    .R0_clk(mem_233_0_R0_clk),
    .R0_data(mem_233_0_R0_data),
    .R0_en(mem_233_0_R0_en),
    .W0_addr(mem_233_0_W0_addr),
    .W0_clk(mem_233_0_W0_clk),
    .W0_data(mem_233_0_W0_data),
    .W0_en(mem_233_0_W0_en),
    .W0_mask(mem_233_0_W0_mask)
  );
  split_mem_0_ext mem_233_1 (
    .R0_addr(mem_233_1_R0_addr),
    .R0_clk(mem_233_1_R0_clk),
    .R0_data(mem_233_1_R0_data),
    .R0_en(mem_233_1_R0_en),
    .W0_addr(mem_233_1_W0_addr),
    .W0_clk(mem_233_1_W0_clk),
    .W0_data(mem_233_1_W0_data),
    .W0_en(mem_233_1_W0_en),
    .W0_mask(mem_233_1_W0_mask)
  );
  split_mem_0_ext mem_233_2 (
    .R0_addr(mem_233_2_R0_addr),
    .R0_clk(mem_233_2_R0_clk),
    .R0_data(mem_233_2_R0_data),
    .R0_en(mem_233_2_R0_en),
    .W0_addr(mem_233_2_W0_addr),
    .W0_clk(mem_233_2_W0_clk),
    .W0_data(mem_233_2_W0_data),
    .W0_en(mem_233_2_W0_en),
    .W0_mask(mem_233_2_W0_mask)
  );
  split_mem_0_ext mem_233_3 (
    .R0_addr(mem_233_3_R0_addr),
    .R0_clk(mem_233_3_R0_clk),
    .R0_data(mem_233_3_R0_data),
    .R0_en(mem_233_3_R0_en),
    .W0_addr(mem_233_3_W0_addr),
    .W0_clk(mem_233_3_W0_clk),
    .W0_data(mem_233_3_W0_data),
    .W0_en(mem_233_3_W0_en),
    .W0_mask(mem_233_3_W0_mask)
  );
  split_mem_0_ext mem_233_4 (
    .R0_addr(mem_233_4_R0_addr),
    .R0_clk(mem_233_4_R0_clk),
    .R0_data(mem_233_4_R0_data),
    .R0_en(mem_233_4_R0_en),
    .W0_addr(mem_233_4_W0_addr),
    .W0_clk(mem_233_4_W0_clk),
    .W0_data(mem_233_4_W0_data),
    .W0_en(mem_233_4_W0_en),
    .W0_mask(mem_233_4_W0_mask)
  );
  split_mem_0_ext mem_233_5 (
    .R0_addr(mem_233_5_R0_addr),
    .R0_clk(mem_233_5_R0_clk),
    .R0_data(mem_233_5_R0_data),
    .R0_en(mem_233_5_R0_en),
    .W0_addr(mem_233_5_W0_addr),
    .W0_clk(mem_233_5_W0_clk),
    .W0_data(mem_233_5_W0_data),
    .W0_en(mem_233_5_W0_en),
    .W0_mask(mem_233_5_W0_mask)
  );
  split_mem_0_ext mem_233_6 (
    .R0_addr(mem_233_6_R0_addr),
    .R0_clk(mem_233_6_R0_clk),
    .R0_data(mem_233_6_R0_data),
    .R0_en(mem_233_6_R0_en),
    .W0_addr(mem_233_6_W0_addr),
    .W0_clk(mem_233_6_W0_clk),
    .W0_data(mem_233_6_W0_data),
    .W0_en(mem_233_6_W0_en),
    .W0_mask(mem_233_6_W0_mask)
  );
  split_mem_0_ext mem_233_7 (
    .R0_addr(mem_233_7_R0_addr),
    .R0_clk(mem_233_7_R0_clk),
    .R0_data(mem_233_7_R0_data),
    .R0_en(mem_233_7_R0_en),
    .W0_addr(mem_233_7_W0_addr),
    .W0_clk(mem_233_7_W0_clk),
    .W0_data(mem_233_7_W0_data),
    .W0_en(mem_233_7_W0_en),
    .W0_mask(mem_233_7_W0_mask)
  );
  split_mem_0_ext mem_234_0 (
    .R0_addr(mem_234_0_R0_addr),
    .R0_clk(mem_234_0_R0_clk),
    .R0_data(mem_234_0_R0_data),
    .R0_en(mem_234_0_R0_en),
    .W0_addr(mem_234_0_W0_addr),
    .W0_clk(mem_234_0_W0_clk),
    .W0_data(mem_234_0_W0_data),
    .W0_en(mem_234_0_W0_en),
    .W0_mask(mem_234_0_W0_mask)
  );
  split_mem_0_ext mem_234_1 (
    .R0_addr(mem_234_1_R0_addr),
    .R0_clk(mem_234_1_R0_clk),
    .R0_data(mem_234_1_R0_data),
    .R0_en(mem_234_1_R0_en),
    .W0_addr(mem_234_1_W0_addr),
    .W0_clk(mem_234_1_W0_clk),
    .W0_data(mem_234_1_W0_data),
    .W0_en(mem_234_1_W0_en),
    .W0_mask(mem_234_1_W0_mask)
  );
  split_mem_0_ext mem_234_2 (
    .R0_addr(mem_234_2_R0_addr),
    .R0_clk(mem_234_2_R0_clk),
    .R0_data(mem_234_2_R0_data),
    .R0_en(mem_234_2_R0_en),
    .W0_addr(mem_234_2_W0_addr),
    .W0_clk(mem_234_2_W0_clk),
    .W0_data(mem_234_2_W0_data),
    .W0_en(mem_234_2_W0_en),
    .W0_mask(mem_234_2_W0_mask)
  );
  split_mem_0_ext mem_234_3 (
    .R0_addr(mem_234_3_R0_addr),
    .R0_clk(mem_234_3_R0_clk),
    .R0_data(mem_234_3_R0_data),
    .R0_en(mem_234_3_R0_en),
    .W0_addr(mem_234_3_W0_addr),
    .W0_clk(mem_234_3_W0_clk),
    .W0_data(mem_234_3_W0_data),
    .W0_en(mem_234_3_W0_en),
    .W0_mask(mem_234_3_W0_mask)
  );
  split_mem_0_ext mem_234_4 (
    .R0_addr(mem_234_4_R0_addr),
    .R0_clk(mem_234_4_R0_clk),
    .R0_data(mem_234_4_R0_data),
    .R0_en(mem_234_4_R0_en),
    .W0_addr(mem_234_4_W0_addr),
    .W0_clk(mem_234_4_W0_clk),
    .W0_data(mem_234_4_W0_data),
    .W0_en(mem_234_4_W0_en),
    .W0_mask(mem_234_4_W0_mask)
  );
  split_mem_0_ext mem_234_5 (
    .R0_addr(mem_234_5_R0_addr),
    .R0_clk(mem_234_5_R0_clk),
    .R0_data(mem_234_5_R0_data),
    .R0_en(mem_234_5_R0_en),
    .W0_addr(mem_234_5_W0_addr),
    .W0_clk(mem_234_5_W0_clk),
    .W0_data(mem_234_5_W0_data),
    .W0_en(mem_234_5_W0_en),
    .W0_mask(mem_234_5_W0_mask)
  );
  split_mem_0_ext mem_234_6 (
    .R0_addr(mem_234_6_R0_addr),
    .R0_clk(mem_234_6_R0_clk),
    .R0_data(mem_234_6_R0_data),
    .R0_en(mem_234_6_R0_en),
    .W0_addr(mem_234_6_W0_addr),
    .W0_clk(mem_234_6_W0_clk),
    .W0_data(mem_234_6_W0_data),
    .W0_en(mem_234_6_W0_en),
    .W0_mask(mem_234_6_W0_mask)
  );
  split_mem_0_ext mem_234_7 (
    .R0_addr(mem_234_7_R0_addr),
    .R0_clk(mem_234_7_R0_clk),
    .R0_data(mem_234_7_R0_data),
    .R0_en(mem_234_7_R0_en),
    .W0_addr(mem_234_7_W0_addr),
    .W0_clk(mem_234_7_W0_clk),
    .W0_data(mem_234_7_W0_data),
    .W0_en(mem_234_7_W0_en),
    .W0_mask(mem_234_7_W0_mask)
  );
  split_mem_0_ext mem_235_0 (
    .R0_addr(mem_235_0_R0_addr),
    .R0_clk(mem_235_0_R0_clk),
    .R0_data(mem_235_0_R0_data),
    .R0_en(mem_235_0_R0_en),
    .W0_addr(mem_235_0_W0_addr),
    .W0_clk(mem_235_0_W0_clk),
    .W0_data(mem_235_0_W0_data),
    .W0_en(mem_235_0_W0_en),
    .W0_mask(mem_235_0_W0_mask)
  );
  split_mem_0_ext mem_235_1 (
    .R0_addr(mem_235_1_R0_addr),
    .R0_clk(mem_235_1_R0_clk),
    .R0_data(mem_235_1_R0_data),
    .R0_en(mem_235_1_R0_en),
    .W0_addr(mem_235_1_W0_addr),
    .W0_clk(mem_235_1_W0_clk),
    .W0_data(mem_235_1_W0_data),
    .W0_en(mem_235_1_W0_en),
    .W0_mask(mem_235_1_W0_mask)
  );
  split_mem_0_ext mem_235_2 (
    .R0_addr(mem_235_2_R0_addr),
    .R0_clk(mem_235_2_R0_clk),
    .R0_data(mem_235_2_R0_data),
    .R0_en(mem_235_2_R0_en),
    .W0_addr(mem_235_2_W0_addr),
    .W0_clk(mem_235_2_W0_clk),
    .W0_data(mem_235_2_W0_data),
    .W0_en(mem_235_2_W0_en),
    .W0_mask(mem_235_2_W0_mask)
  );
  split_mem_0_ext mem_235_3 (
    .R0_addr(mem_235_3_R0_addr),
    .R0_clk(mem_235_3_R0_clk),
    .R0_data(mem_235_3_R0_data),
    .R0_en(mem_235_3_R0_en),
    .W0_addr(mem_235_3_W0_addr),
    .W0_clk(mem_235_3_W0_clk),
    .W0_data(mem_235_3_W0_data),
    .W0_en(mem_235_3_W0_en),
    .W0_mask(mem_235_3_W0_mask)
  );
  split_mem_0_ext mem_235_4 (
    .R0_addr(mem_235_4_R0_addr),
    .R0_clk(mem_235_4_R0_clk),
    .R0_data(mem_235_4_R0_data),
    .R0_en(mem_235_4_R0_en),
    .W0_addr(mem_235_4_W0_addr),
    .W0_clk(mem_235_4_W0_clk),
    .W0_data(mem_235_4_W0_data),
    .W0_en(mem_235_4_W0_en),
    .W0_mask(mem_235_4_W0_mask)
  );
  split_mem_0_ext mem_235_5 (
    .R0_addr(mem_235_5_R0_addr),
    .R0_clk(mem_235_5_R0_clk),
    .R0_data(mem_235_5_R0_data),
    .R0_en(mem_235_5_R0_en),
    .W0_addr(mem_235_5_W0_addr),
    .W0_clk(mem_235_5_W0_clk),
    .W0_data(mem_235_5_W0_data),
    .W0_en(mem_235_5_W0_en),
    .W0_mask(mem_235_5_W0_mask)
  );
  split_mem_0_ext mem_235_6 (
    .R0_addr(mem_235_6_R0_addr),
    .R0_clk(mem_235_6_R0_clk),
    .R0_data(mem_235_6_R0_data),
    .R0_en(mem_235_6_R0_en),
    .W0_addr(mem_235_6_W0_addr),
    .W0_clk(mem_235_6_W0_clk),
    .W0_data(mem_235_6_W0_data),
    .W0_en(mem_235_6_W0_en),
    .W0_mask(mem_235_6_W0_mask)
  );
  split_mem_0_ext mem_235_7 (
    .R0_addr(mem_235_7_R0_addr),
    .R0_clk(mem_235_7_R0_clk),
    .R0_data(mem_235_7_R0_data),
    .R0_en(mem_235_7_R0_en),
    .W0_addr(mem_235_7_W0_addr),
    .W0_clk(mem_235_7_W0_clk),
    .W0_data(mem_235_7_W0_data),
    .W0_en(mem_235_7_W0_en),
    .W0_mask(mem_235_7_W0_mask)
  );
  split_mem_0_ext mem_236_0 (
    .R0_addr(mem_236_0_R0_addr),
    .R0_clk(mem_236_0_R0_clk),
    .R0_data(mem_236_0_R0_data),
    .R0_en(mem_236_0_R0_en),
    .W0_addr(mem_236_0_W0_addr),
    .W0_clk(mem_236_0_W0_clk),
    .W0_data(mem_236_0_W0_data),
    .W0_en(mem_236_0_W0_en),
    .W0_mask(mem_236_0_W0_mask)
  );
  split_mem_0_ext mem_236_1 (
    .R0_addr(mem_236_1_R0_addr),
    .R0_clk(mem_236_1_R0_clk),
    .R0_data(mem_236_1_R0_data),
    .R0_en(mem_236_1_R0_en),
    .W0_addr(mem_236_1_W0_addr),
    .W0_clk(mem_236_1_W0_clk),
    .W0_data(mem_236_1_W0_data),
    .W0_en(mem_236_1_W0_en),
    .W0_mask(mem_236_1_W0_mask)
  );
  split_mem_0_ext mem_236_2 (
    .R0_addr(mem_236_2_R0_addr),
    .R0_clk(mem_236_2_R0_clk),
    .R0_data(mem_236_2_R0_data),
    .R0_en(mem_236_2_R0_en),
    .W0_addr(mem_236_2_W0_addr),
    .W0_clk(mem_236_2_W0_clk),
    .W0_data(mem_236_2_W0_data),
    .W0_en(mem_236_2_W0_en),
    .W0_mask(mem_236_2_W0_mask)
  );
  split_mem_0_ext mem_236_3 (
    .R0_addr(mem_236_3_R0_addr),
    .R0_clk(mem_236_3_R0_clk),
    .R0_data(mem_236_3_R0_data),
    .R0_en(mem_236_3_R0_en),
    .W0_addr(mem_236_3_W0_addr),
    .W0_clk(mem_236_3_W0_clk),
    .W0_data(mem_236_3_W0_data),
    .W0_en(mem_236_3_W0_en),
    .W0_mask(mem_236_3_W0_mask)
  );
  split_mem_0_ext mem_236_4 (
    .R0_addr(mem_236_4_R0_addr),
    .R0_clk(mem_236_4_R0_clk),
    .R0_data(mem_236_4_R0_data),
    .R0_en(mem_236_4_R0_en),
    .W0_addr(mem_236_4_W0_addr),
    .W0_clk(mem_236_4_W0_clk),
    .W0_data(mem_236_4_W0_data),
    .W0_en(mem_236_4_W0_en),
    .W0_mask(mem_236_4_W0_mask)
  );
  split_mem_0_ext mem_236_5 (
    .R0_addr(mem_236_5_R0_addr),
    .R0_clk(mem_236_5_R0_clk),
    .R0_data(mem_236_5_R0_data),
    .R0_en(mem_236_5_R0_en),
    .W0_addr(mem_236_5_W0_addr),
    .W0_clk(mem_236_5_W0_clk),
    .W0_data(mem_236_5_W0_data),
    .W0_en(mem_236_5_W0_en),
    .W0_mask(mem_236_5_W0_mask)
  );
  split_mem_0_ext mem_236_6 (
    .R0_addr(mem_236_6_R0_addr),
    .R0_clk(mem_236_6_R0_clk),
    .R0_data(mem_236_6_R0_data),
    .R0_en(mem_236_6_R0_en),
    .W0_addr(mem_236_6_W0_addr),
    .W0_clk(mem_236_6_W0_clk),
    .W0_data(mem_236_6_W0_data),
    .W0_en(mem_236_6_W0_en),
    .W0_mask(mem_236_6_W0_mask)
  );
  split_mem_0_ext mem_236_7 (
    .R0_addr(mem_236_7_R0_addr),
    .R0_clk(mem_236_7_R0_clk),
    .R0_data(mem_236_7_R0_data),
    .R0_en(mem_236_7_R0_en),
    .W0_addr(mem_236_7_W0_addr),
    .W0_clk(mem_236_7_W0_clk),
    .W0_data(mem_236_7_W0_data),
    .W0_en(mem_236_7_W0_en),
    .W0_mask(mem_236_7_W0_mask)
  );
  split_mem_0_ext mem_237_0 (
    .R0_addr(mem_237_0_R0_addr),
    .R0_clk(mem_237_0_R0_clk),
    .R0_data(mem_237_0_R0_data),
    .R0_en(mem_237_0_R0_en),
    .W0_addr(mem_237_0_W0_addr),
    .W0_clk(mem_237_0_W0_clk),
    .W0_data(mem_237_0_W0_data),
    .W0_en(mem_237_0_W0_en),
    .W0_mask(mem_237_0_W0_mask)
  );
  split_mem_0_ext mem_237_1 (
    .R0_addr(mem_237_1_R0_addr),
    .R0_clk(mem_237_1_R0_clk),
    .R0_data(mem_237_1_R0_data),
    .R0_en(mem_237_1_R0_en),
    .W0_addr(mem_237_1_W0_addr),
    .W0_clk(mem_237_1_W0_clk),
    .W0_data(mem_237_1_W0_data),
    .W0_en(mem_237_1_W0_en),
    .W0_mask(mem_237_1_W0_mask)
  );
  split_mem_0_ext mem_237_2 (
    .R0_addr(mem_237_2_R0_addr),
    .R0_clk(mem_237_2_R0_clk),
    .R0_data(mem_237_2_R0_data),
    .R0_en(mem_237_2_R0_en),
    .W0_addr(mem_237_2_W0_addr),
    .W0_clk(mem_237_2_W0_clk),
    .W0_data(mem_237_2_W0_data),
    .W0_en(mem_237_2_W0_en),
    .W0_mask(mem_237_2_W0_mask)
  );
  split_mem_0_ext mem_237_3 (
    .R0_addr(mem_237_3_R0_addr),
    .R0_clk(mem_237_3_R0_clk),
    .R0_data(mem_237_3_R0_data),
    .R0_en(mem_237_3_R0_en),
    .W0_addr(mem_237_3_W0_addr),
    .W0_clk(mem_237_3_W0_clk),
    .W0_data(mem_237_3_W0_data),
    .W0_en(mem_237_3_W0_en),
    .W0_mask(mem_237_3_W0_mask)
  );
  split_mem_0_ext mem_237_4 (
    .R0_addr(mem_237_4_R0_addr),
    .R0_clk(mem_237_4_R0_clk),
    .R0_data(mem_237_4_R0_data),
    .R0_en(mem_237_4_R0_en),
    .W0_addr(mem_237_4_W0_addr),
    .W0_clk(mem_237_4_W0_clk),
    .W0_data(mem_237_4_W0_data),
    .W0_en(mem_237_4_W0_en),
    .W0_mask(mem_237_4_W0_mask)
  );
  split_mem_0_ext mem_237_5 (
    .R0_addr(mem_237_5_R0_addr),
    .R0_clk(mem_237_5_R0_clk),
    .R0_data(mem_237_5_R0_data),
    .R0_en(mem_237_5_R0_en),
    .W0_addr(mem_237_5_W0_addr),
    .W0_clk(mem_237_5_W0_clk),
    .W0_data(mem_237_5_W0_data),
    .W0_en(mem_237_5_W0_en),
    .W0_mask(mem_237_5_W0_mask)
  );
  split_mem_0_ext mem_237_6 (
    .R0_addr(mem_237_6_R0_addr),
    .R0_clk(mem_237_6_R0_clk),
    .R0_data(mem_237_6_R0_data),
    .R0_en(mem_237_6_R0_en),
    .W0_addr(mem_237_6_W0_addr),
    .W0_clk(mem_237_6_W0_clk),
    .W0_data(mem_237_6_W0_data),
    .W0_en(mem_237_6_W0_en),
    .W0_mask(mem_237_6_W0_mask)
  );
  split_mem_0_ext mem_237_7 (
    .R0_addr(mem_237_7_R0_addr),
    .R0_clk(mem_237_7_R0_clk),
    .R0_data(mem_237_7_R0_data),
    .R0_en(mem_237_7_R0_en),
    .W0_addr(mem_237_7_W0_addr),
    .W0_clk(mem_237_7_W0_clk),
    .W0_data(mem_237_7_W0_data),
    .W0_en(mem_237_7_W0_en),
    .W0_mask(mem_237_7_W0_mask)
  );
  split_mem_0_ext mem_238_0 (
    .R0_addr(mem_238_0_R0_addr),
    .R0_clk(mem_238_0_R0_clk),
    .R0_data(mem_238_0_R0_data),
    .R0_en(mem_238_0_R0_en),
    .W0_addr(mem_238_0_W0_addr),
    .W0_clk(mem_238_0_W0_clk),
    .W0_data(mem_238_0_W0_data),
    .W0_en(mem_238_0_W0_en),
    .W0_mask(mem_238_0_W0_mask)
  );
  split_mem_0_ext mem_238_1 (
    .R0_addr(mem_238_1_R0_addr),
    .R0_clk(mem_238_1_R0_clk),
    .R0_data(mem_238_1_R0_data),
    .R0_en(mem_238_1_R0_en),
    .W0_addr(mem_238_1_W0_addr),
    .W0_clk(mem_238_1_W0_clk),
    .W0_data(mem_238_1_W0_data),
    .W0_en(mem_238_1_W0_en),
    .W0_mask(mem_238_1_W0_mask)
  );
  split_mem_0_ext mem_238_2 (
    .R0_addr(mem_238_2_R0_addr),
    .R0_clk(mem_238_2_R0_clk),
    .R0_data(mem_238_2_R0_data),
    .R0_en(mem_238_2_R0_en),
    .W0_addr(mem_238_2_W0_addr),
    .W0_clk(mem_238_2_W0_clk),
    .W0_data(mem_238_2_W0_data),
    .W0_en(mem_238_2_W0_en),
    .W0_mask(mem_238_2_W0_mask)
  );
  split_mem_0_ext mem_238_3 (
    .R0_addr(mem_238_3_R0_addr),
    .R0_clk(mem_238_3_R0_clk),
    .R0_data(mem_238_3_R0_data),
    .R0_en(mem_238_3_R0_en),
    .W0_addr(mem_238_3_W0_addr),
    .W0_clk(mem_238_3_W0_clk),
    .W0_data(mem_238_3_W0_data),
    .W0_en(mem_238_3_W0_en),
    .W0_mask(mem_238_3_W0_mask)
  );
  split_mem_0_ext mem_238_4 (
    .R0_addr(mem_238_4_R0_addr),
    .R0_clk(mem_238_4_R0_clk),
    .R0_data(mem_238_4_R0_data),
    .R0_en(mem_238_4_R0_en),
    .W0_addr(mem_238_4_W0_addr),
    .W0_clk(mem_238_4_W0_clk),
    .W0_data(mem_238_4_W0_data),
    .W0_en(mem_238_4_W0_en),
    .W0_mask(mem_238_4_W0_mask)
  );
  split_mem_0_ext mem_238_5 (
    .R0_addr(mem_238_5_R0_addr),
    .R0_clk(mem_238_5_R0_clk),
    .R0_data(mem_238_5_R0_data),
    .R0_en(mem_238_5_R0_en),
    .W0_addr(mem_238_5_W0_addr),
    .W0_clk(mem_238_5_W0_clk),
    .W0_data(mem_238_5_W0_data),
    .W0_en(mem_238_5_W0_en),
    .W0_mask(mem_238_5_W0_mask)
  );
  split_mem_0_ext mem_238_6 (
    .R0_addr(mem_238_6_R0_addr),
    .R0_clk(mem_238_6_R0_clk),
    .R0_data(mem_238_6_R0_data),
    .R0_en(mem_238_6_R0_en),
    .W0_addr(mem_238_6_W0_addr),
    .W0_clk(mem_238_6_W0_clk),
    .W0_data(mem_238_6_W0_data),
    .W0_en(mem_238_6_W0_en),
    .W0_mask(mem_238_6_W0_mask)
  );
  split_mem_0_ext mem_238_7 (
    .R0_addr(mem_238_7_R0_addr),
    .R0_clk(mem_238_7_R0_clk),
    .R0_data(mem_238_7_R0_data),
    .R0_en(mem_238_7_R0_en),
    .W0_addr(mem_238_7_W0_addr),
    .W0_clk(mem_238_7_W0_clk),
    .W0_data(mem_238_7_W0_data),
    .W0_en(mem_238_7_W0_en),
    .W0_mask(mem_238_7_W0_mask)
  );
  split_mem_0_ext mem_239_0 (
    .R0_addr(mem_239_0_R0_addr),
    .R0_clk(mem_239_0_R0_clk),
    .R0_data(mem_239_0_R0_data),
    .R0_en(mem_239_0_R0_en),
    .W0_addr(mem_239_0_W0_addr),
    .W0_clk(mem_239_0_W0_clk),
    .W0_data(mem_239_0_W0_data),
    .W0_en(mem_239_0_W0_en),
    .W0_mask(mem_239_0_W0_mask)
  );
  split_mem_0_ext mem_239_1 (
    .R0_addr(mem_239_1_R0_addr),
    .R0_clk(mem_239_1_R0_clk),
    .R0_data(mem_239_1_R0_data),
    .R0_en(mem_239_1_R0_en),
    .W0_addr(mem_239_1_W0_addr),
    .W0_clk(mem_239_1_W0_clk),
    .W0_data(mem_239_1_W0_data),
    .W0_en(mem_239_1_W0_en),
    .W0_mask(mem_239_1_W0_mask)
  );
  split_mem_0_ext mem_239_2 (
    .R0_addr(mem_239_2_R0_addr),
    .R0_clk(mem_239_2_R0_clk),
    .R0_data(mem_239_2_R0_data),
    .R0_en(mem_239_2_R0_en),
    .W0_addr(mem_239_2_W0_addr),
    .W0_clk(mem_239_2_W0_clk),
    .W0_data(mem_239_2_W0_data),
    .W0_en(mem_239_2_W0_en),
    .W0_mask(mem_239_2_W0_mask)
  );
  split_mem_0_ext mem_239_3 (
    .R0_addr(mem_239_3_R0_addr),
    .R0_clk(mem_239_3_R0_clk),
    .R0_data(mem_239_3_R0_data),
    .R0_en(mem_239_3_R0_en),
    .W0_addr(mem_239_3_W0_addr),
    .W0_clk(mem_239_3_W0_clk),
    .W0_data(mem_239_3_W0_data),
    .W0_en(mem_239_3_W0_en),
    .W0_mask(mem_239_3_W0_mask)
  );
  split_mem_0_ext mem_239_4 (
    .R0_addr(mem_239_4_R0_addr),
    .R0_clk(mem_239_4_R0_clk),
    .R0_data(mem_239_4_R0_data),
    .R0_en(mem_239_4_R0_en),
    .W0_addr(mem_239_4_W0_addr),
    .W0_clk(mem_239_4_W0_clk),
    .W0_data(mem_239_4_W0_data),
    .W0_en(mem_239_4_W0_en),
    .W0_mask(mem_239_4_W0_mask)
  );
  split_mem_0_ext mem_239_5 (
    .R0_addr(mem_239_5_R0_addr),
    .R0_clk(mem_239_5_R0_clk),
    .R0_data(mem_239_5_R0_data),
    .R0_en(mem_239_5_R0_en),
    .W0_addr(mem_239_5_W0_addr),
    .W0_clk(mem_239_5_W0_clk),
    .W0_data(mem_239_5_W0_data),
    .W0_en(mem_239_5_W0_en),
    .W0_mask(mem_239_5_W0_mask)
  );
  split_mem_0_ext mem_239_6 (
    .R0_addr(mem_239_6_R0_addr),
    .R0_clk(mem_239_6_R0_clk),
    .R0_data(mem_239_6_R0_data),
    .R0_en(mem_239_6_R0_en),
    .W0_addr(mem_239_6_W0_addr),
    .W0_clk(mem_239_6_W0_clk),
    .W0_data(mem_239_6_W0_data),
    .W0_en(mem_239_6_W0_en),
    .W0_mask(mem_239_6_W0_mask)
  );
  split_mem_0_ext mem_239_7 (
    .R0_addr(mem_239_7_R0_addr),
    .R0_clk(mem_239_7_R0_clk),
    .R0_data(mem_239_7_R0_data),
    .R0_en(mem_239_7_R0_en),
    .W0_addr(mem_239_7_W0_addr),
    .W0_clk(mem_239_7_W0_clk),
    .W0_data(mem_239_7_W0_data),
    .W0_en(mem_239_7_W0_en),
    .W0_mask(mem_239_7_W0_mask)
  );
  split_mem_0_ext mem_240_0 (
    .R0_addr(mem_240_0_R0_addr),
    .R0_clk(mem_240_0_R0_clk),
    .R0_data(mem_240_0_R0_data),
    .R0_en(mem_240_0_R0_en),
    .W0_addr(mem_240_0_W0_addr),
    .W0_clk(mem_240_0_W0_clk),
    .W0_data(mem_240_0_W0_data),
    .W0_en(mem_240_0_W0_en),
    .W0_mask(mem_240_0_W0_mask)
  );
  split_mem_0_ext mem_240_1 (
    .R0_addr(mem_240_1_R0_addr),
    .R0_clk(mem_240_1_R0_clk),
    .R0_data(mem_240_1_R0_data),
    .R0_en(mem_240_1_R0_en),
    .W0_addr(mem_240_1_W0_addr),
    .W0_clk(mem_240_1_W0_clk),
    .W0_data(mem_240_1_W0_data),
    .W0_en(mem_240_1_W0_en),
    .W0_mask(mem_240_1_W0_mask)
  );
  split_mem_0_ext mem_240_2 (
    .R0_addr(mem_240_2_R0_addr),
    .R0_clk(mem_240_2_R0_clk),
    .R0_data(mem_240_2_R0_data),
    .R0_en(mem_240_2_R0_en),
    .W0_addr(mem_240_2_W0_addr),
    .W0_clk(mem_240_2_W0_clk),
    .W0_data(mem_240_2_W0_data),
    .W0_en(mem_240_2_W0_en),
    .W0_mask(mem_240_2_W0_mask)
  );
  split_mem_0_ext mem_240_3 (
    .R0_addr(mem_240_3_R0_addr),
    .R0_clk(mem_240_3_R0_clk),
    .R0_data(mem_240_3_R0_data),
    .R0_en(mem_240_3_R0_en),
    .W0_addr(mem_240_3_W0_addr),
    .W0_clk(mem_240_3_W0_clk),
    .W0_data(mem_240_3_W0_data),
    .W0_en(mem_240_3_W0_en),
    .W0_mask(mem_240_3_W0_mask)
  );
  split_mem_0_ext mem_240_4 (
    .R0_addr(mem_240_4_R0_addr),
    .R0_clk(mem_240_4_R0_clk),
    .R0_data(mem_240_4_R0_data),
    .R0_en(mem_240_4_R0_en),
    .W0_addr(mem_240_4_W0_addr),
    .W0_clk(mem_240_4_W0_clk),
    .W0_data(mem_240_4_W0_data),
    .W0_en(mem_240_4_W0_en),
    .W0_mask(mem_240_4_W0_mask)
  );
  split_mem_0_ext mem_240_5 (
    .R0_addr(mem_240_5_R0_addr),
    .R0_clk(mem_240_5_R0_clk),
    .R0_data(mem_240_5_R0_data),
    .R0_en(mem_240_5_R0_en),
    .W0_addr(mem_240_5_W0_addr),
    .W0_clk(mem_240_5_W0_clk),
    .W0_data(mem_240_5_W0_data),
    .W0_en(mem_240_5_W0_en),
    .W0_mask(mem_240_5_W0_mask)
  );
  split_mem_0_ext mem_240_6 (
    .R0_addr(mem_240_6_R0_addr),
    .R0_clk(mem_240_6_R0_clk),
    .R0_data(mem_240_6_R0_data),
    .R0_en(mem_240_6_R0_en),
    .W0_addr(mem_240_6_W0_addr),
    .W0_clk(mem_240_6_W0_clk),
    .W0_data(mem_240_6_W0_data),
    .W0_en(mem_240_6_W0_en),
    .W0_mask(mem_240_6_W0_mask)
  );
  split_mem_0_ext mem_240_7 (
    .R0_addr(mem_240_7_R0_addr),
    .R0_clk(mem_240_7_R0_clk),
    .R0_data(mem_240_7_R0_data),
    .R0_en(mem_240_7_R0_en),
    .W0_addr(mem_240_7_W0_addr),
    .W0_clk(mem_240_7_W0_clk),
    .W0_data(mem_240_7_W0_data),
    .W0_en(mem_240_7_W0_en),
    .W0_mask(mem_240_7_W0_mask)
  );
  split_mem_0_ext mem_241_0 (
    .R0_addr(mem_241_0_R0_addr),
    .R0_clk(mem_241_0_R0_clk),
    .R0_data(mem_241_0_R0_data),
    .R0_en(mem_241_0_R0_en),
    .W0_addr(mem_241_0_W0_addr),
    .W0_clk(mem_241_0_W0_clk),
    .W0_data(mem_241_0_W0_data),
    .W0_en(mem_241_0_W0_en),
    .W0_mask(mem_241_0_W0_mask)
  );
  split_mem_0_ext mem_241_1 (
    .R0_addr(mem_241_1_R0_addr),
    .R0_clk(mem_241_1_R0_clk),
    .R0_data(mem_241_1_R0_data),
    .R0_en(mem_241_1_R0_en),
    .W0_addr(mem_241_1_W0_addr),
    .W0_clk(mem_241_1_W0_clk),
    .W0_data(mem_241_1_W0_data),
    .W0_en(mem_241_1_W0_en),
    .W0_mask(mem_241_1_W0_mask)
  );
  split_mem_0_ext mem_241_2 (
    .R0_addr(mem_241_2_R0_addr),
    .R0_clk(mem_241_2_R0_clk),
    .R0_data(mem_241_2_R0_data),
    .R0_en(mem_241_2_R0_en),
    .W0_addr(mem_241_2_W0_addr),
    .W0_clk(mem_241_2_W0_clk),
    .W0_data(mem_241_2_W0_data),
    .W0_en(mem_241_2_W0_en),
    .W0_mask(mem_241_2_W0_mask)
  );
  split_mem_0_ext mem_241_3 (
    .R0_addr(mem_241_3_R0_addr),
    .R0_clk(mem_241_3_R0_clk),
    .R0_data(mem_241_3_R0_data),
    .R0_en(mem_241_3_R0_en),
    .W0_addr(mem_241_3_W0_addr),
    .W0_clk(mem_241_3_W0_clk),
    .W0_data(mem_241_3_W0_data),
    .W0_en(mem_241_3_W0_en),
    .W0_mask(mem_241_3_W0_mask)
  );
  split_mem_0_ext mem_241_4 (
    .R0_addr(mem_241_4_R0_addr),
    .R0_clk(mem_241_4_R0_clk),
    .R0_data(mem_241_4_R0_data),
    .R0_en(mem_241_4_R0_en),
    .W0_addr(mem_241_4_W0_addr),
    .W0_clk(mem_241_4_W0_clk),
    .W0_data(mem_241_4_W0_data),
    .W0_en(mem_241_4_W0_en),
    .W0_mask(mem_241_4_W0_mask)
  );
  split_mem_0_ext mem_241_5 (
    .R0_addr(mem_241_5_R0_addr),
    .R0_clk(mem_241_5_R0_clk),
    .R0_data(mem_241_5_R0_data),
    .R0_en(mem_241_5_R0_en),
    .W0_addr(mem_241_5_W0_addr),
    .W0_clk(mem_241_5_W0_clk),
    .W0_data(mem_241_5_W0_data),
    .W0_en(mem_241_5_W0_en),
    .W0_mask(mem_241_5_W0_mask)
  );
  split_mem_0_ext mem_241_6 (
    .R0_addr(mem_241_6_R0_addr),
    .R0_clk(mem_241_6_R0_clk),
    .R0_data(mem_241_6_R0_data),
    .R0_en(mem_241_6_R0_en),
    .W0_addr(mem_241_6_W0_addr),
    .W0_clk(mem_241_6_W0_clk),
    .W0_data(mem_241_6_W0_data),
    .W0_en(mem_241_6_W0_en),
    .W0_mask(mem_241_6_W0_mask)
  );
  split_mem_0_ext mem_241_7 (
    .R0_addr(mem_241_7_R0_addr),
    .R0_clk(mem_241_7_R0_clk),
    .R0_data(mem_241_7_R0_data),
    .R0_en(mem_241_7_R0_en),
    .W0_addr(mem_241_7_W0_addr),
    .W0_clk(mem_241_7_W0_clk),
    .W0_data(mem_241_7_W0_data),
    .W0_en(mem_241_7_W0_en),
    .W0_mask(mem_241_7_W0_mask)
  );
  split_mem_0_ext mem_242_0 (
    .R0_addr(mem_242_0_R0_addr),
    .R0_clk(mem_242_0_R0_clk),
    .R0_data(mem_242_0_R0_data),
    .R0_en(mem_242_0_R0_en),
    .W0_addr(mem_242_0_W0_addr),
    .W0_clk(mem_242_0_W0_clk),
    .W0_data(mem_242_0_W0_data),
    .W0_en(mem_242_0_W0_en),
    .W0_mask(mem_242_0_W0_mask)
  );
  split_mem_0_ext mem_242_1 (
    .R0_addr(mem_242_1_R0_addr),
    .R0_clk(mem_242_1_R0_clk),
    .R0_data(mem_242_1_R0_data),
    .R0_en(mem_242_1_R0_en),
    .W0_addr(mem_242_1_W0_addr),
    .W0_clk(mem_242_1_W0_clk),
    .W0_data(mem_242_1_W0_data),
    .W0_en(mem_242_1_W0_en),
    .W0_mask(mem_242_1_W0_mask)
  );
  split_mem_0_ext mem_242_2 (
    .R0_addr(mem_242_2_R0_addr),
    .R0_clk(mem_242_2_R0_clk),
    .R0_data(mem_242_2_R0_data),
    .R0_en(mem_242_2_R0_en),
    .W0_addr(mem_242_2_W0_addr),
    .W0_clk(mem_242_2_W0_clk),
    .W0_data(mem_242_2_W0_data),
    .W0_en(mem_242_2_W0_en),
    .W0_mask(mem_242_2_W0_mask)
  );
  split_mem_0_ext mem_242_3 (
    .R0_addr(mem_242_3_R0_addr),
    .R0_clk(mem_242_3_R0_clk),
    .R0_data(mem_242_3_R0_data),
    .R0_en(mem_242_3_R0_en),
    .W0_addr(mem_242_3_W0_addr),
    .W0_clk(mem_242_3_W0_clk),
    .W0_data(mem_242_3_W0_data),
    .W0_en(mem_242_3_W0_en),
    .W0_mask(mem_242_3_W0_mask)
  );
  split_mem_0_ext mem_242_4 (
    .R0_addr(mem_242_4_R0_addr),
    .R0_clk(mem_242_4_R0_clk),
    .R0_data(mem_242_4_R0_data),
    .R0_en(mem_242_4_R0_en),
    .W0_addr(mem_242_4_W0_addr),
    .W0_clk(mem_242_4_W0_clk),
    .W0_data(mem_242_4_W0_data),
    .W0_en(mem_242_4_W0_en),
    .W0_mask(mem_242_4_W0_mask)
  );
  split_mem_0_ext mem_242_5 (
    .R0_addr(mem_242_5_R0_addr),
    .R0_clk(mem_242_5_R0_clk),
    .R0_data(mem_242_5_R0_data),
    .R0_en(mem_242_5_R0_en),
    .W0_addr(mem_242_5_W0_addr),
    .W0_clk(mem_242_5_W0_clk),
    .W0_data(mem_242_5_W0_data),
    .W0_en(mem_242_5_W0_en),
    .W0_mask(mem_242_5_W0_mask)
  );
  split_mem_0_ext mem_242_6 (
    .R0_addr(mem_242_6_R0_addr),
    .R0_clk(mem_242_6_R0_clk),
    .R0_data(mem_242_6_R0_data),
    .R0_en(mem_242_6_R0_en),
    .W0_addr(mem_242_6_W0_addr),
    .W0_clk(mem_242_6_W0_clk),
    .W0_data(mem_242_6_W0_data),
    .W0_en(mem_242_6_W0_en),
    .W0_mask(mem_242_6_W0_mask)
  );
  split_mem_0_ext mem_242_7 (
    .R0_addr(mem_242_7_R0_addr),
    .R0_clk(mem_242_7_R0_clk),
    .R0_data(mem_242_7_R0_data),
    .R0_en(mem_242_7_R0_en),
    .W0_addr(mem_242_7_W0_addr),
    .W0_clk(mem_242_7_W0_clk),
    .W0_data(mem_242_7_W0_data),
    .W0_en(mem_242_7_W0_en),
    .W0_mask(mem_242_7_W0_mask)
  );
  split_mem_0_ext mem_243_0 (
    .R0_addr(mem_243_0_R0_addr),
    .R0_clk(mem_243_0_R0_clk),
    .R0_data(mem_243_0_R0_data),
    .R0_en(mem_243_0_R0_en),
    .W0_addr(mem_243_0_W0_addr),
    .W0_clk(mem_243_0_W0_clk),
    .W0_data(mem_243_0_W0_data),
    .W0_en(mem_243_0_W0_en),
    .W0_mask(mem_243_0_W0_mask)
  );
  split_mem_0_ext mem_243_1 (
    .R0_addr(mem_243_1_R0_addr),
    .R0_clk(mem_243_1_R0_clk),
    .R0_data(mem_243_1_R0_data),
    .R0_en(mem_243_1_R0_en),
    .W0_addr(mem_243_1_W0_addr),
    .W0_clk(mem_243_1_W0_clk),
    .W0_data(mem_243_1_W0_data),
    .W0_en(mem_243_1_W0_en),
    .W0_mask(mem_243_1_W0_mask)
  );
  split_mem_0_ext mem_243_2 (
    .R0_addr(mem_243_2_R0_addr),
    .R0_clk(mem_243_2_R0_clk),
    .R0_data(mem_243_2_R0_data),
    .R0_en(mem_243_2_R0_en),
    .W0_addr(mem_243_2_W0_addr),
    .W0_clk(mem_243_2_W0_clk),
    .W0_data(mem_243_2_W0_data),
    .W0_en(mem_243_2_W0_en),
    .W0_mask(mem_243_2_W0_mask)
  );
  split_mem_0_ext mem_243_3 (
    .R0_addr(mem_243_3_R0_addr),
    .R0_clk(mem_243_3_R0_clk),
    .R0_data(mem_243_3_R0_data),
    .R0_en(mem_243_3_R0_en),
    .W0_addr(mem_243_3_W0_addr),
    .W0_clk(mem_243_3_W0_clk),
    .W0_data(mem_243_3_W0_data),
    .W0_en(mem_243_3_W0_en),
    .W0_mask(mem_243_3_W0_mask)
  );
  split_mem_0_ext mem_243_4 (
    .R0_addr(mem_243_4_R0_addr),
    .R0_clk(mem_243_4_R0_clk),
    .R0_data(mem_243_4_R0_data),
    .R0_en(mem_243_4_R0_en),
    .W0_addr(mem_243_4_W0_addr),
    .W0_clk(mem_243_4_W0_clk),
    .W0_data(mem_243_4_W0_data),
    .W0_en(mem_243_4_W0_en),
    .W0_mask(mem_243_4_W0_mask)
  );
  split_mem_0_ext mem_243_5 (
    .R0_addr(mem_243_5_R0_addr),
    .R0_clk(mem_243_5_R0_clk),
    .R0_data(mem_243_5_R0_data),
    .R0_en(mem_243_5_R0_en),
    .W0_addr(mem_243_5_W0_addr),
    .W0_clk(mem_243_5_W0_clk),
    .W0_data(mem_243_5_W0_data),
    .W0_en(mem_243_5_W0_en),
    .W0_mask(mem_243_5_W0_mask)
  );
  split_mem_0_ext mem_243_6 (
    .R0_addr(mem_243_6_R0_addr),
    .R0_clk(mem_243_6_R0_clk),
    .R0_data(mem_243_6_R0_data),
    .R0_en(mem_243_6_R0_en),
    .W0_addr(mem_243_6_W0_addr),
    .W0_clk(mem_243_6_W0_clk),
    .W0_data(mem_243_6_W0_data),
    .W0_en(mem_243_6_W0_en),
    .W0_mask(mem_243_6_W0_mask)
  );
  split_mem_0_ext mem_243_7 (
    .R0_addr(mem_243_7_R0_addr),
    .R0_clk(mem_243_7_R0_clk),
    .R0_data(mem_243_7_R0_data),
    .R0_en(mem_243_7_R0_en),
    .W0_addr(mem_243_7_W0_addr),
    .W0_clk(mem_243_7_W0_clk),
    .W0_data(mem_243_7_W0_data),
    .W0_en(mem_243_7_W0_en),
    .W0_mask(mem_243_7_W0_mask)
  );
  split_mem_0_ext mem_244_0 (
    .R0_addr(mem_244_0_R0_addr),
    .R0_clk(mem_244_0_R0_clk),
    .R0_data(mem_244_0_R0_data),
    .R0_en(mem_244_0_R0_en),
    .W0_addr(mem_244_0_W0_addr),
    .W0_clk(mem_244_0_W0_clk),
    .W0_data(mem_244_0_W0_data),
    .W0_en(mem_244_0_W0_en),
    .W0_mask(mem_244_0_W0_mask)
  );
  split_mem_0_ext mem_244_1 (
    .R0_addr(mem_244_1_R0_addr),
    .R0_clk(mem_244_1_R0_clk),
    .R0_data(mem_244_1_R0_data),
    .R0_en(mem_244_1_R0_en),
    .W0_addr(mem_244_1_W0_addr),
    .W0_clk(mem_244_1_W0_clk),
    .W0_data(mem_244_1_W0_data),
    .W0_en(mem_244_1_W0_en),
    .W0_mask(mem_244_1_W0_mask)
  );
  split_mem_0_ext mem_244_2 (
    .R0_addr(mem_244_2_R0_addr),
    .R0_clk(mem_244_2_R0_clk),
    .R0_data(mem_244_2_R0_data),
    .R0_en(mem_244_2_R0_en),
    .W0_addr(mem_244_2_W0_addr),
    .W0_clk(mem_244_2_W0_clk),
    .W0_data(mem_244_2_W0_data),
    .W0_en(mem_244_2_W0_en),
    .W0_mask(mem_244_2_W0_mask)
  );
  split_mem_0_ext mem_244_3 (
    .R0_addr(mem_244_3_R0_addr),
    .R0_clk(mem_244_3_R0_clk),
    .R0_data(mem_244_3_R0_data),
    .R0_en(mem_244_3_R0_en),
    .W0_addr(mem_244_3_W0_addr),
    .W0_clk(mem_244_3_W0_clk),
    .W0_data(mem_244_3_W0_data),
    .W0_en(mem_244_3_W0_en),
    .W0_mask(mem_244_3_W0_mask)
  );
  split_mem_0_ext mem_244_4 (
    .R0_addr(mem_244_4_R0_addr),
    .R0_clk(mem_244_4_R0_clk),
    .R0_data(mem_244_4_R0_data),
    .R0_en(mem_244_4_R0_en),
    .W0_addr(mem_244_4_W0_addr),
    .W0_clk(mem_244_4_W0_clk),
    .W0_data(mem_244_4_W0_data),
    .W0_en(mem_244_4_W0_en),
    .W0_mask(mem_244_4_W0_mask)
  );
  split_mem_0_ext mem_244_5 (
    .R0_addr(mem_244_5_R0_addr),
    .R0_clk(mem_244_5_R0_clk),
    .R0_data(mem_244_5_R0_data),
    .R0_en(mem_244_5_R0_en),
    .W0_addr(mem_244_5_W0_addr),
    .W0_clk(mem_244_5_W0_clk),
    .W0_data(mem_244_5_W0_data),
    .W0_en(mem_244_5_W0_en),
    .W0_mask(mem_244_5_W0_mask)
  );
  split_mem_0_ext mem_244_6 (
    .R0_addr(mem_244_6_R0_addr),
    .R0_clk(mem_244_6_R0_clk),
    .R0_data(mem_244_6_R0_data),
    .R0_en(mem_244_6_R0_en),
    .W0_addr(mem_244_6_W0_addr),
    .W0_clk(mem_244_6_W0_clk),
    .W0_data(mem_244_6_W0_data),
    .W0_en(mem_244_6_W0_en),
    .W0_mask(mem_244_6_W0_mask)
  );
  split_mem_0_ext mem_244_7 (
    .R0_addr(mem_244_7_R0_addr),
    .R0_clk(mem_244_7_R0_clk),
    .R0_data(mem_244_7_R0_data),
    .R0_en(mem_244_7_R0_en),
    .W0_addr(mem_244_7_W0_addr),
    .W0_clk(mem_244_7_W0_clk),
    .W0_data(mem_244_7_W0_data),
    .W0_en(mem_244_7_W0_en),
    .W0_mask(mem_244_7_W0_mask)
  );
  split_mem_0_ext mem_245_0 (
    .R0_addr(mem_245_0_R0_addr),
    .R0_clk(mem_245_0_R0_clk),
    .R0_data(mem_245_0_R0_data),
    .R0_en(mem_245_0_R0_en),
    .W0_addr(mem_245_0_W0_addr),
    .W0_clk(mem_245_0_W0_clk),
    .W0_data(mem_245_0_W0_data),
    .W0_en(mem_245_0_W0_en),
    .W0_mask(mem_245_0_W0_mask)
  );
  split_mem_0_ext mem_245_1 (
    .R0_addr(mem_245_1_R0_addr),
    .R0_clk(mem_245_1_R0_clk),
    .R0_data(mem_245_1_R0_data),
    .R0_en(mem_245_1_R0_en),
    .W0_addr(mem_245_1_W0_addr),
    .W0_clk(mem_245_1_W0_clk),
    .W0_data(mem_245_1_W0_data),
    .W0_en(mem_245_1_W0_en),
    .W0_mask(mem_245_1_W0_mask)
  );
  split_mem_0_ext mem_245_2 (
    .R0_addr(mem_245_2_R0_addr),
    .R0_clk(mem_245_2_R0_clk),
    .R0_data(mem_245_2_R0_data),
    .R0_en(mem_245_2_R0_en),
    .W0_addr(mem_245_2_W0_addr),
    .W0_clk(mem_245_2_W0_clk),
    .W0_data(mem_245_2_W0_data),
    .W0_en(mem_245_2_W0_en),
    .W0_mask(mem_245_2_W0_mask)
  );
  split_mem_0_ext mem_245_3 (
    .R0_addr(mem_245_3_R0_addr),
    .R0_clk(mem_245_3_R0_clk),
    .R0_data(mem_245_3_R0_data),
    .R0_en(mem_245_3_R0_en),
    .W0_addr(mem_245_3_W0_addr),
    .W0_clk(mem_245_3_W0_clk),
    .W0_data(mem_245_3_W0_data),
    .W0_en(mem_245_3_W0_en),
    .W0_mask(mem_245_3_W0_mask)
  );
  split_mem_0_ext mem_245_4 (
    .R0_addr(mem_245_4_R0_addr),
    .R0_clk(mem_245_4_R0_clk),
    .R0_data(mem_245_4_R0_data),
    .R0_en(mem_245_4_R0_en),
    .W0_addr(mem_245_4_W0_addr),
    .W0_clk(mem_245_4_W0_clk),
    .W0_data(mem_245_4_W0_data),
    .W0_en(mem_245_4_W0_en),
    .W0_mask(mem_245_4_W0_mask)
  );
  split_mem_0_ext mem_245_5 (
    .R0_addr(mem_245_5_R0_addr),
    .R0_clk(mem_245_5_R0_clk),
    .R0_data(mem_245_5_R0_data),
    .R0_en(mem_245_5_R0_en),
    .W0_addr(mem_245_5_W0_addr),
    .W0_clk(mem_245_5_W0_clk),
    .W0_data(mem_245_5_W0_data),
    .W0_en(mem_245_5_W0_en),
    .W0_mask(mem_245_5_W0_mask)
  );
  split_mem_0_ext mem_245_6 (
    .R0_addr(mem_245_6_R0_addr),
    .R0_clk(mem_245_6_R0_clk),
    .R0_data(mem_245_6_R0_data),
    .R0_en(mem_245_6_R0_en),
    .W0_addr(mem_245_6_W0_addr),
    .W0_clk(mem_245_6_W0_clk),
    .W0_data(mem_245_6_W0_data),
    .W0_en(mem_245_6_W0_en),
    .W0_mask(mem_245_6_W0_mask)
  );
  split_mem_0_ext mem_245_7 (
    .R0_addr(mem_245_7_R0_addr),
    .R0_clk(mem_245_7_R0_clk),
    .R0_data(mem_245_7_R0_data),
    .R0_en(mem_245_7_R0_en),
    .W0_addr(mem_245_7_W0_addr),
    .W0_clk(mem_245_7_W0_clk),
    .W0_data(mem_245_7_W0_data),
    .W0_en(mem_245_7_W0_en),
    .W0_mask(mem_245_7_W0_mask)
  );
  split_mem_0_ext mem_246_0 (
    .R0_addr(mem_246_0_R0_addr),
    .R0_clk(mem_246_0_R0_clk),
    .R0_data(mem_246_0_R0_data),
    .R0_en(mem_246_0_R0_en),
    .W0_addr(mem_246_0_W0_addr),
    .W0_clk(mem_246_0_W0_clk),
    .W0_data(mem_246_0_W0_data),
    .W0_en(mem_246_0_W0_en),
    .W0_mask(mem_246_0_W0_mask)
  );
  split_mem_0_ext mem_246_1 (
    .R0_addr(mem_246_1_R0_addr),
    .R0_clk(mem_246_1_R0_clk),
    .R0_data(mem_246_1_R0_data),
    .R0_en(mem_246_1_R0_en),
    .W0_addr(mem_246_1_W0_addr),
    .W0_clk(mem_246_1_W0_clk),
    .W0_data(mem_246_1_W0_data),
    .W0_en(mem_246_1_W0_en),
    .W0_mask(mem_246_1_W0_mask)
  );
  split_mem_0_ext mem_246_2 (
    .R0_addr(mem_246_2_R0_addr),
    .R0_clk(mem_246_2_R0_clk),
    .R0_data(mem_246_2_R0_data),
    .R0_en(mem_246_2_R0_en),
    .W0_addr(mem_246_2_W0_addr),
    .W0_clk(mem_246_2_W0_clk),
    .W0_data(mem_246_2_W0_data),
    .W0_en(mem_246_2_W0_en),
    .W0_mask(mem_246_2_W0_mask)
  );
  split_mem_0_ext mem_246_3 (
    .R0_addr(mem_246_3_R0_addr),
    .R0_clk(mem_246_3_R0_clk),
    .R0_data(mem_246_3_R0_data),
    .R0_en(mem_246_3_R0_en),
    .W0_addr(mem_246_3_W0_addr),
    .W0_clk(mem_246_3_W0_clk),
    .W0_data(mem_246_3_W0_data),
    .W0_en(mem_246_3_W0_en),
    .W0_mask(mem_246_3_W0_mask)
  );
  split_mem_0_ext mem_246_4 (
    .R0_addr(mem_246_4_R0_addr),
    .R0_clk(mem_246_4_R0_clk),
    .R0_data(mem_246_4_R0_data),
    .R0_en(mem_246_4_R0_en),
    .W0_addr(mem_246_4_W0_addr),
    .W0_clk(mem_246_4_W0_clk),
    .W0_data(mem_246_4_W0_data),
    .W0_en(mem_246_4_W0_en),
    .W0_mask(mem_246_4_W0_mask)
  );
  split_mem_0_ext mem_246_5 (
    .R0_addr(mem_246_5_R0_addr),
    .R0_clk(mem_246_5_R0_clk),
    .R0_data(mem_246_5_R0_data),
    .R0_en(mem_246_5_R0_en),
    .W0_addr(mem_246_5_W0_addr),
    .W0_clk(mem_246_5_W0_clk),
    .W0_data(mem_246_5_W0_data),
    .W0_en(mem_246_5_W0_en),
    .W0_mask(mem_246_5_W0_mask)
  );
  split_mem_0_ext mem_246_6 (
    .R0_addr(mem_246_6_R0_addr),
    .R0_clk(mem_246_6_R0_clk),
    .R0_data(mem_246_6_R0_data),
    .R0_en(mem_246_6_R0_en),
    .W0_addr(mem_246_6_W0_addr),
    .W0_clk(mem_246_6_W0_clk),
    .W0_data(mem_246_6_W0_data),
    .W0_en(mem_246_6_W0_en),
    .W0_mask(mem_246_6_W0_mask)
  );
  split_mem_0_ext mem_246_7 (
    .R0_addr(mem_246_7_R0_addr),
    .R0_clk(mem_246_7_R0_clk),
    .R0_data(mem_246_7_R0_data),
    .R0_en(mem_246_7_R0_en),
    .W0_addr(mem_246_7_W0_addr),
    .W0_clk(mem_246_7_W0_clk),
    .W0_data(mem_246_7_W0_data),
    .W0_en(mem_246_7_W0_en),
    .W0_mask(mem_246_7_W0_mask)
  );
  split_mem_0_ext mem_247_0 (
    .R0_addr(mem_247_0_R0_addr),
    .R0_clk(mem_247_0_R0_clk),
    .R0_data(mem_247_0_R0_data),
    .R0_en(mem_247_0_R0_en),
    .W0_addr(mem_247_0_W0_addr),
    .W0_clk(mem_247_0_W0_clk),
    .W0_data(mem_247_0_W0_data),
    .W0_en(mem_247_0_W0_en),
    .W0_mask(mem_247_0_W0_mask)
  );
  split_mem_0_ext mem_247_1 (
    .R0_addr(mem_247_1_R0_addr),
    .R0_clk(mem_247_1_R0_clk),
    .R0_data(mem_247_1_R0_data),
    .R0_en(mem_247_1_R0_en),
    .W0_addr(mem_247_1_W0_addr),
    .W0_clk(mem_247_1_W0_clk),
    .W0_data(mem_247_1_W0_data),
    .W0_en(mem_247_1_W0_en),
    .W0_mask(mem_247_1_W0_mask)
  );
  split_mem_0_ext mem_247_2 (
    .R0_addr(mem_247_2_R0_addr),
    .R0_clk(mem_247_2_R0_clk),
    .R0_data(mem_247_2_R0_data),
    .R0_en(mem_247_2_R0_en),
    .W0_addr(mem_247_2_W0_addr),
    .W0_clk(mem_247_2_W0_clk),
    .W0_data(mem_247_2_W0_data),
    .W0_en(mem_247_2_W0_en),
    .W0_mask(mem_247_2_W0_mask)
  );
  split_mem_0_ext mem_247_3 (
    .R0_addr(mem_247_3_R0_addr),
    .R0_clk(mem_247_3_R0_clk),
    .R0_data(mem_247_3_R0_data),
    .R0_en(mem_247_3_R0_en),
    .W0_addr(mem_247_3_W0_addr),
    .W0_clk(mem_247_3_W0_clk),
    .W0_data(mem_247_3_W0_data),
    .W0_en(mem_247_3_W0_en),
    .W0_mask(mem_247_3_W0_mask)
  );
  split_mem_0_ext mem_247_4 (
    .R0_addr(mem_247_4_R0_addr),
    .R0_clk(mem_247_4_R0_clk),
    .R0_data(mem_247_4_R0_data),
    .R0_en(mem_247_4_R0_en),
    .W0_addr(mem_247_4_W0_addr),
    .W0_clk(mem_247_4_W0_clk),
    .W0_data(mem_247_4_W0_data),
    .W0_en(mem_247_4_W0_en),
    .W0_mask(mem_247_4_W0_mask)
  );
  split_mem_0_ext mem_247_5 (
    .R0_addr(mem_247_5_R0_addr),
    .R0_clk(mem_247_5_R0_clk),
    .R0_data(mem_247_5_R0_data),
    .R0_en(mem_247_5_R0_en),
    .W0_addr(mem_247_5_W0_addr),
    .W0_clk(mem_247_5_W0_clk),
    .W0_data(mem_247_5_W0_data),
    .W0_en(mem_247_5_W0_en),
    .W0_mask(mem_247_5_W0_mask)
  );
  split_mem_0_ext mem_247_6 (
    .R0_addr(mem_247_6_R0_addr),
    .R0_clk(mem_247_6_R0_clk),
    .R0_data(mem_247_6_R0_data),
    .R0_en(mem_247_6_R0_en),
    .W0_addr(mem_247_6_W0_addr),
    .W0_clk(mem_247_6_W0_clk),
    .W0_data(mem_247_6_W0_data),
    .W0_en(mem_247_6_W0_en),
    .W0_mask(mem_247_6_W0_mask)
  );
  split_mem_0_ext mem_247_7 (
    .R0_addr(mem_247_7_R0_addr),
    .R0_clk(mem_247_7_R0_clk),
    .R0_data(mem_247_7_R0_data),
    .R0_en(mem_247_7_R0_en),
    .W0_addr(mem_247_7_W0_addr),
    .W0_clk(mem_247_7_W0_clk),
    .W0_data(mem_247_7_W0_data),
    .W0_en(mem_247_7_W0_en),
    .W0_mask(mem_247_7_W0_mask)
  );
  split_mem_0_ext mem_248_0 (
    .R0_addr(mem_248_0_R0_addr),
    .R0_clk(mem_248_0_R0_clk),
    .R0_data(mem_248_0_R0_data),
    .R0_en(mem_248_0_R0_en),
    .W0_addr(mem_248_0_W0_addr),
    .W0_clk(mem_248_0_W0_clk),
    .W0_data(mem_248_0_W0_data),
    .W0_en(mem_248_0_W0_en),
    .W0_mask(mem_248_0_W0_mask)
  );
  split_mem_0_ext mem_248_1 (
    .R0_addr(mem_248_1_R0_addr),
    .R0_clk(mem_248_1_R0_clk),
    .R0_data(mem_248_1_R0_data),
    .R0_en(mem_248_1_R0_en),
    .W0_addr(mem_248_1_W0_addr),
    .W0_clk(mem_248_1_W0_clk),
    .W0_data(mem_248_1_W0_data),
    .W0_en(mem_248_1_W0_en),
    .W0_mask(mem_248_1_W0_mask)
  );
  split_mem_0_ext mem_248_2 (
    .R0_addr(mem_248_2_R0_addr),
    .R0_clk(mem_248_2_R0_clk),
    .R0_data(mem_248_2_R0_data),
    .R0_en(mem_248_2_R0_en),
    .W0_addr(mem_248_2_W0_addr),
    .W0_clk(mem_248_2_W0_clk),
    .W0_data(mem_248_2_W0_data),
    .W0_en(mem_248_2_W0_en),
    .W0_mask(mem_248_2_W0_mask)
  );
  split_mem_0_ext mem_248_3 (
    .R0_addr(mem_248_3_R0_addr),
    .R0_clk(mem_248_3_R0_clk),
    .R0_data(mem_248_3_R0_data),
    .R0_en(mem_248_3_R0_en),
    .W0_addr(mem_248_3_W0_addr),
    .W0_clk(mem_248_3_W0_clk),
    .W0_data(mem_248_3_W0_data),
    .W0_en(mem_248_3_W0_en),
    .W0_mask(mem_248_3_W0_mask)
  );
  split_mem_0_ext mem_248_4 (
    .R0_addr(mem_248_4_R0_addr),
    .R0_clk(mem_248_4_R0_clk),
    .R0_data(mem_248_4_R0_data),
    .R0_en(mem_248_4_R0_en),
    .W0_addr(mem_248_4_W0_addr),
    .W0_clk(mem_248_4_W0_clk),
    .W0_data(mem_248_4_W0_data),
    .W0_en(mem_248_4_W0_en),
    .W0_mask(mem_248_4_W0_mask)
  );
  split_mem_0_ext mem_248_5 (
    .R0_addr(mem_248_5_R0_addr),
    .R0_clk(mem_248_5_R0_clk),
    .R0_data(mem_248_5_R0_data),
    .R0_en(mem_248_5_R0_en),
    .W0_addr(mem_248_5_W0_addr),
    .W0_clk(mem_248_5_W0_clk),
    .W0_data(mem_248_5_W0_data),
    .W0_en(mem_248_5_W0_en),
    .W0_mask(mem_248_5_W0_mask)
  );
  split_mem_0_ext mem_248_6 (
    .R0_addr(mem_248_6_R0_addr),
    .R0_clk(mem_248_6_R0_clk),
    .R0_data(mem_248_6_R0_data),
    .R0_en(mem_248_6_R0_en),
    .W0_addr(mem_248_6_W0_addr),
    .W0_clk(mem_248_6_W0_clk),
    .W0_data(mem_248_6_W0_data),
    .W0_en(mem_248_6_W0_en),
    .W0_mask(mem_248_6_W0_mask)
  );
  split_mem_0_ext mem_248_7 (
    .R0_addr(mem_248_7_R0_addr),
    .R0_clk(mem_248_7_R0_clk),
    .R0_data(mem_248_7_R0_data),
    .R0_en(mem_248_7_R0_en),
    .W0_addr(mem_248_7_W0_addr),
    .W0_clk(mem_248_7_W0_clk),
    .W0_data(mem_248_7_W0_data),
    .W0_en(mem_248_7_W0_en),
    .W0_mask(mem_248_7_W0_mask)
  );
  split_mem_0_ext mem_249_0 (
    .R0_addr(mem_249_0_R0_addr),
    .R0_clk(mem_249_0_R0_clk),
    .R0_data(mem_249_0_R0_data),
    .R0_en(mem_249_0_R0_en),
    .W0_addr(mem_249_0_W0_addr),
    .W0_clk(mem_249_0_W0_clk),
    .W0_data(mem_249_0_W0_data),
    .W0_en(mem_249_0_W0_en),
    .W0_mask(mem_249_0_W0_mask)
  );
  split_mem_0_ext mem_249_1 (
    .R0_addr(mem_249_1_R0_addr),
    .R0_clk(mem_249_1_R0_clk),
    .R0_data(mem_249_1_R0_data),
    .R0_en(mem_249_1_R0_en),
    .W0_addr(mem_249_1_W0_addr),
    .W0_clk(mem_249_1_W0_clk),
    .W0_data(mem_249_1_W0_data),
    .W0_en(mem_249_1_W0_en),
    .W0_mask(mem_249_1_W0_mask)
  );
  split_mem_0_ext mem_249_2 (
    .R0_addr(mem_249_2_R0_addr),
    .R0_clk(mem_249_2_R0_clk),
    .R0_data(mem_249_2_R0_data),
    .R0_en(mem_249_2_R0_en),
    .W0_addr(mem_249_2_W0_addr),
    .W0_clk(mem_249_2_W0_clk),
    .W0_data(mem_249_2_W0_data),
    .W0_en(mem_249_2_W0_en),
    .W0_mask(mem_249_2_W0_mask)
  );
  split_mem_0_ext mem_249_3 (
    .R0_addr(mem_249_3_R0_addr),
    .R0_clk(mem_249_3_R0_clk),
    .R0_data(mem_249_3_R0_data),
    .R0_en(mem_249_3_R0_en),
    .W0_addr(mem_249_3_W0_addr),
    .W0_clk(mem_249_3_W0_clk),
    .W0_data(mem_249_3_W0_data),
    .W0_en(mem_249_3_W0_en),
    .W0_mask(mem_249_3_W0_mask)
  );
  split_mem_0_ext mem_249_4 (
    .R0_addr(mem_249_4_R0_addr),
    .R0_clk(mem_249_4_R0_clk),
    .R0_data(mem_249_4_R0_data),
    .R0_en(mem_249_4_R0_en),
    .W0_addr(mem_249_4_W0_addr),
    .W0_clk(mem_249_4_W0_clk),
    .W0_data(mem_249_4_W0_data),
    .W0_en(mem_249_4_W0_en),
    .W0_mask(mem_249_4_W0_mask)
  );
  split_mem_0_ext mem_249_5 (
    .R0_addr(mem_249_5_R0_addr),
    .R0_clk(mem_249_5_R0_clk),
    .R0_data(mem_249_5_R0_data),
    .R0_en(mem_249_5_R0_en),
    .W0_addr(mem_249_5_W0_addr),
    .W0_clk(mem_249_5_W0_clk),
    .W0_data(mem_249_5_W0_data),
    .W0_en(mem_249_5_W0_en),
    .W0_mask(mem_249_5_W0_mask)
  );
  split_mem_0_ext mem_249_6 (
    .R0_addr(mem_249_6_R0_addr),
    .R0_clk(mem_249_6_R0_clk),
    .R0_data(mem_249_6_R0_data),
    .R0_en(mem_249_6_R0_en),
    .W0_addr(mem_249_6_W0_addr),
    .W0_clk(mem_249_6_W0_clk),
    .W0_data(mem_249_6_W0_data),
    .W0_en(mem_249_6_W0_en),
    .W0_mask(mem_249_6_W0_mask)
  );
  split_mem_0_ext mem_249_7 (
    .R0_addr(mem_249_7_R0_addr),
    .R0_clk(mem_249_7_R0_clk),
    .R0_data(mem_249_7_R0_data),
    .R0_en(mem_249_7_R0_en),
    .W0_addr(mem_249_7_W0_addr),
    .W0_clk(mem_249_7_W0_clk),
    .W0_data(mem_249_7_W0_data),
    .W0_en(mem_249_7_W0_en),
    .W0_mask(mem_249_7_W0_mask)
  );
  split_mem_0_ext mem_250_0 (
    .R0_addr(mem_250_0_R0_addr),
    .R0_clk(mem_250_0_R0_clk),
    .R0_data(mem_250_0_R0_data),
    .R0_en(mem_250_0_R0_en),
    .W0_addr(mem_250_0_W0_addr),
    .W0_clk(mem_250_0_W0_clk),
    .W0_data(mem_250_0_W0_data),
    .W0_en(mem_250_0_W0_en),
    .W0_mask(mem_250_0_W0_mask)
  );
  split_mem_0_ext mem_250_1 (
    .R0_addr(mem_250_1_R0_addr),
    .R0_clk(mem_250_1_R0_clk),
    .R0_data(mem_250_1_R0_data),
    .R0_en(mem_250_1_R0_en),
    .W0_addr(mem_250_1_W0_addr),
    .W0_clk(mem_250_1_W0_clk),
    .W0_data(mem_250_1_W0_data),
    .W0_en(mem_250_1_W0_en),
    .W0_mask(mem_250_1_W0_mask)
  );
  split_mem_0_ext mem_250_2 (
    .R0_addr(mem_250_2_R0_addr),
    .R0_clk(mem_250_2_R0_clk),
    .R0_data(mem_250_2_R0_data),
    .R0_en(mem_250_2_R0_en),
    .W0_addr(mem_250_2_W0_addr),
    .W0_clk(mem_250_2_W0_clk),
    .W0_data(mem_250_2_W0_data),
    .W0_en(mem_250_2_W0_en),
    .W0_mask(mem_250_2_W0_mask)
  );
  split_mem_0_ext mem_250_3 (
    .R0_addr(mem_250_3_R0_addr),
    .R0_clk(mem_250_3_R0_clk),
    .R0_data(mem_250_3_R0_data),
    .R0_en(mem_250_3_R0_en),
    .W0_addr(mem_250_3_W0_addr),
    .W0_clk(mem_250_3_W0_clk),
    .W0_data(mem_250_3_W0_data),
    .W0_en(mem_250_3_W0_en),
    .W0_mask(mem_250_3_W0_mask)
  );
  split_mem_0_ext mem_250_4 (
    .R0_addr(mem_250_4_R0_addr),
    .R0_clk(mem_250_4_R0_clk),
    .R0_data(mem_250_4_R0_data),
    .R0_en(mem_250_4_R0_en),
    .W0_addr(mem_250_4_W0_addr),
    .W0_clk(mem_250_4_W0_clk),
    .W0_data(mem_250_4_W0_data),
    .W0_en(mem_250_4_W0_en),
    .W0_mask(mem_250_4_W0_mask)
  );
  split_mem_0_ext mem_250_5 (
    .R0_addr(mem_250_5_R0_addr),
    .R0_clk(mem_250_5_R0_clk),
    .R0_data(mem_250_5_R0_data),
    .R0_en(mem_250_5_R0_en),
    .W0_addr(mem_250_5_W0_addr),
    .W0_clk(mem_250_5_W0_clk),
    .W0_data(mem_250_5_W0_data),
    .W0_en(mem_250_5_W0_en),
    .W0_mask(mem_250_5_W0_mask)
  );
  split_mem_0_ext mem_250_6 (
    .R0_addr(mem_250_6_R0_addr),
    .R0_clk(mem_250_6_R0_clk),
    .R0_data(mem_250_6_R0_data),
    .R0_en(mem_250_6_R0_en),
    .W0_addr(mem_250_6_W0_addr),
    .W0_clk(mem_250_6_W0_clk),
    .W0_data(mem_250_6_W0_data),
    .W0_en(mem_250_6_W0_en),
    .W0_mask(mem_250_6_W0_mask)
  );
  split_mem_0_ext mem_250_7 (
    .R0_addr(mem_250_7_R0_addr),
    .R0_clk(mem_250_7_R0_clk),
    .R0_data(mem_250_7_R0_data),
    .R0_en(mem_250_7_R0_en),
    .W0_addr(mem_250_7_W0_addr),
    .W0_clk(mem_250_7_W0_clk),
    .W0_data(mem_250_7_W0_data),
    .W0_en(mem_250_7_W0_en),
    .W0_mask(mem_250_7_W0_mask)
  );
  split_mem_0_ext mem_251_0 (
    .R0_addr(mem_251_0_R0_addr),
    .R0_clk(mem_251_0_R0_clk),
    .R0_data(mem_251_0_R0_data),
    .R0_en(mem_251_0_R0_en),
    .W0_addr(mem_251_0_W0_addr),
    .W0_clk(mem_251_0_W0_clk),
    .W0_data(mem_251_0_W0_data),
    .W0_en(mem_251_0_W0_en),
    .W0_mask(mem_251_0_W0_mask)
  );
  split_mem_0_ext mem_251_1 (
    .R0_addr(mem_251_1_R0_addr),
    .R0_clk(mem_251_1_R0_clk),
    .R0_data(mem_251_1_R0_data),
    .R0_en(mem_251_1_R0_en),
    .W0_addr(mem_251_1_W0_addr),
    .W0_clk(mem_251_1_W0_clk),
    .W0_data(mem_251_1_W0_data),
    .W0_en(mem_251_1_W0_en),
    .W0_mask(mem_251_1_W0_mask)
  );
  split_mem_0_ext mem_251_2 (
    .R0_addr(mem_251_2_R0_addr),
    .R0_clk(mem_251_2_R0_clk),
    .R0_data(mem_251_2_R0_data),
    .R0_en(mem_251_2_R0_en),
    .W0_addr(mem_251_2_W0_addr),
    .W0_clk(mem_251_2_W0_clk),
    .W0_data(mem_251_2_W0_data),
    .W0_en(mem_251_2_W0_en),
    .W0_mask(mem_251_2_W0_mask)
  );
  split_mem_0_ext mem_251_3 (
    .R0_addr(mem_251_3_R0_addr),
    .R0_clk(mem_251_3_R0_clk),
    .R0_data(mem_251_3_R0_data),
    .R0_en(mem_251_3_R0_en),
    .W0_addr(mem_251_3_W0_addr),
    .W0_clk(mem_251_3_W0_clk),
    .W0_data(mem_251_3_W0_data),
    .W0_en(mem_251_3_W0_en),
    .W0_mask(mem_251_3_W0_mask)
  );
  split_mem_0_ext mem_251_4 (
    .R0_addr(mem_251_4_R0_addr),
    .R0_clk(mem_251_4_R0_clk),
    .R0_data(mem_251_4_R0_data),
    .R0_en(mem_251_4_R0_en),
    .W0_addr(mem_251_4_W0_addr),
    .W0_clk(mem_251_4_W0_clk),
    .W0_data(mem_251_4_W0_data),
    .W0_en(mem_251_4_W0_en),
    .W0_mask(mem_251_4_W0_mask)
  );
  split_mem_0_ext mem_251_5 (
    .R0_addr(mem_251_5_R0_addr),
    .R0_clk(mem_251_5_R0_clk),
    .R0_data(mem_251_5_R0_data),
    .R0_en(mem_251_5_R0_en),
    .W0_addr(mem_251_5_W0_addr),
    .W0_clk(mem_251_5_W0_clk),
    .W0_data(mem_251_5_W0_data),
    .W0_en(mem_251_5_W0_en),
    .W0_mask(mem_251_5_W0_mask)
  );
  split_mem_0_ext mem_251_6 (
    .R0_addr(mem_251_6_R0_addr),
    .R0_clk(mem_251_6_R0_clk),
    .R0_data(mem_251_6_R0_data),
    .R0_en(mem_251_6_R0_en),
    .W0_addr(mem_251_6_W0_addr),
    .W0_clk(mem_251_6_W0_clk),
    .W0_data(mem_251_6_W0_data),
    .W0_en(mem_251_6_W0_en),
    .W0_mask(mem_251_6_W0_mask)
  );
  split_mem_0_ext mem_251_7 (
    .R0_addr(mem_251_7_R0_addr),
    .R0_clk(mem_251_7_R0_clk),
    .R0_data(mem_251_7_R0_data),
    .R0_en(mem_251_7_R0_en),
    .W0_addr(mem_251_7_W0_addr),
    .W0_clk(mem_251_7_W0_clk),
    .W0_data(mem_251_7_W0_data),
    .W0_en(mem_251_7_W0_en),
    .W0_mask(mem_251_7_W0_mask)
  );
  split_mem_0_ext mem_252_0 (
    .R0_addr(mem_252_0_R0_addr),
    .R0_clk(mem_252_0_R0_clk),
    .R0_data(mem_252_0_R0_data),
    .R0_en(mem_252_0_R0_en),
    .W0_addr(mem_252_0_W0_addr),
    .W0_clk(mem_252_0_W0_clk),
    .W0_data(mem_252_0_W0_data),
    .W0_en(mem_252_0_W0_en),
    .W0_mask(mem_252_0_W0_mask)
  );
  split_mem_0_ext mem_252_1 (
    .R0_addr(mem_252_1_R0_addr),
    .R0_clk(mem_252_1_R0_clk),
    .R0_data(mem_252_1_R0_data),
    .R0_en(mem_252_1_R0_en),
    .W0_addr(mem_252_1_W0_addr),
    .W0_clk(mem_252_1_W0_clk),
    .W0_data(mem_252_1_W0_data),
    .W0_en(mem_252_1_W0_en),
    .W0_mask(mem_252_1_W0_mask)
  );
  split_mem_0_ext mem_252_2 (
    .R0_addr(mem_252_2_R0_addr),
    .R0_clk(mem_252_2_R0_clk),
    .R0_data(mem_252_2_R0_data),
    .R0_en(mem_252_2_R0_en),
    .W0_addr(mem_252_2_W0_addr),
    .W0_clk(mem_252_2_W0_clk),
    .W0_data(mem_252_2_W0_data),
    .W0_en(mem_252_2_W0_en),
    .W0_mask(mem_252_2_W0_mask)
  );
  split_mem_0_ext mem_252_3 (
    .R0_addr(mem_252_3_R0_addr),
    .R0_clk(mem_252_3_R0_clk),
    .R0_data(mem_252_3_R0_data),
    .R0_en(mem_252_3_R0_en),
    .W0_addr(mem_252_3_W0_addr),
    .W0_clk(mem_252_3_W0_clk),
    .W0_data(mem_252_3_W0_data),
    .W0_en(mem_252_3_W0_en),
    .W0_mask(mem_252_3_W0_mask)
  );
  split_mem_0_ext mem_252_4 (
    .R0_addr(mem_252_4_R0_addr),
    .R0_clk(mem_252_4_R0_clk),
    .R0_data(mem_252_4_R0_data),
    .R0_en(mem_252_4_R0_en),
    .W0_addr(mem_252_4_W0_addr),
    .W0_clk(mem_252_4_W0_clk),
    .W0_data(mem_252_4_W0_data),
    .W0_en(mem_252_4_W0_en),
    .W0_mask(mem_252_4_W0_mask)
  );
  split_mem_0_ext mem_252_5 (
    .R0_addr(mem_252_5_R0_addr),
    .R0_clk(mem_252_5_R0_clk),
    .R0_data(mem_252_5_R0_data),
    .R0_en(mem_252_5_R0_en),
    .W0_addr(mem_252_5_W0_addr),
    .W0_clk(mem_252_5_W0_clk),
    .W0_data(mem_252_5_W0_data),
    .W0_en(mem_252_5_W0_en),
    .W0_mask(mem_252_5_W0_mask)
  );
  split_mem_0_ext mem_252_6 (
    .R0_addr(mem_252_6_R0_addr),
    .R0_clk(mem_252_6_R0_clk),
    .R0_data(mem_252_6_R0_data),
    .R0_en(mem_252_6_R0_en),
    .W0_addr(mem_252_6_W0_addr),
    .W0_clk(mem_252_6_W0_clk),
    .W0_data(mem_252_6_W0_data),
    .W0_en(mem_252_6_W0_en),
    .W0_mask(mem_252_6_W0_mask)
  );
  split_mem_0_ext mem_252_7 (
    .R0_addr(mem_252_7_R0_addr),
    .R0_clk(mem_252_7_R0_clk),
    .R0_data(mem_252_7_R0_data),
    .R0_en(mem_252_7_R0_en),
    .W0_addr(mem_252_7_W0_addr),
    .W0_clk(mem_252_7_W0_clk),
    .W0_data(mem_252_7_W0_data),
    .W0_en(mem_252_7_W0_en),
    .W0_mask(mem_252_7_W0_mask)
  );
  split_mem_0_ext mem_253_0 (
    .R0_addr(mem_253_0_R0_addr),
    .R0_clk(mem_253_0_R0_clk),
    .R0_data(mem_253_0_R0_data),
    .R0_en(mem_253_0_R0_en),
    .W0_addr(mem_253_0_W0_addr),
    .W0_clk(mem_253_0_W0_clk),
    .W0_data(mem_253_0_W0_data),
    .W0_en(mem_253_0_W0_en),
    .W0_mask(mem_253_0_W0_mask)
  );
  split_mem_0_ext mem_253_1 (
    .R0_addr(mem_253_1_R0_addr),
    .R0_clk(mem_253_1_R0_clk),
    .R0_data(mem_253_1_R0_data),
    .R0_en(mem_253_1_R0_en),
    .W0_addr(mem_253_1_W0_addr),
    .W0_clk(mem_253_1_W0_clk),
    .W0_data(mem_253_1_W0_data),
    .W0_en(mem_253_1_W0_en),
    .W0_mask(mem_253_1_W0_mask)
  );
  split_mem_0_ext mem_253_2 (
    .R0_addr(mem_253_2_R0_addr),
    .R0_clk(mem_253_2_R0_clk),
    .R0_data(mem_253_2_R0_data),
    .R0_en(mem_253_2_R0_en),
    .W0_addr(mem_253_2_W0_addr),
    .W0_clk(mem_253_2_W0_clk),
    .W0_data(mem_253_2_W0_data),
    .W0_en(mem_253_2_W0_en),
    .W0_mask(mem_253_2_W0_mask)
  );
  split_mem_0_ext mem_253_3 (
    .R0_addr(mem_253_3_R0_addr),
    .R0_clk(mem_253_3_R0_clk),
    .R0_data(mem_253_3_R0_data),
    .R0_en(mem_253_3_R0_en),
    .W0_addr(mem_253_3_W0_addr),
    .W0_clk(mem_253_3_W0_clk),
    .W0_data(mem_253_3_W0_data),
    .W0_en(mem_253_3_W0_en),
    .W0_mask(mem_253_3_W0_mask)
  );
  split_mem_0_ext mem_253_4 (
    .R0_addr(mem_253_4_R0_addr),
    .R0_clk(mem_253_4_R0_clk),
    .R0_data(mem_253_4_R0_data),
    .R0_en(mem_253_4_R0_en),
    .W0_addr(mem_253_4_W0_addr),
    .W0_clk(mem_253_4_W0_clk),
    .W0_data(mem_253_4_W0_data),
    .W0_en(mem_253_4_W0_en),
    .W0_mask(mem_253_4_W0_mask)
  );
  split_mem_0_ext mem_253_5 (
    .R0_addr(mem_253_5_R0_addr),
    .R0_clk(mem_253_5_R0_clk),
    .R0_data(mem_253_5_R0_data),
    .R0_en(mem_253_5_R0_en),
    .W0_addr(mem_253_5_W0_addr),
    .W0_clk(mem_253_5_W0_clk),
    .W0_data(mem_253_5_W0_data),
    .W0_en(mem_253_5_W0_en),
    .W0_mask(mem_253_5_W0_mask)
  );
  split_mem_0_ext mem_253_6 (
    .R0_addr(mem_253_6_R0_addr),
    .R0_clk(mem_253_6_R0_clk),
    .R0_data(mem_253_6_R0_data),
    .R0_en(mem_253_6_R0_en),
    .W0_addr(mem_253_6_W0_addr),
    .W0_clk(mem_253_6_W0_clk),
    .W0_data(mem_253_6_W0_data),
    .W0_en(mem_253_6_W0_en),
    .W0_mask(mem_253_6_W0_mask)
  );
  split_mem_0_ext mem_253_7 (
    .R0_addr(mem_253_7_R0_addr),
    .R0_clk(mem_253_7_R0_clk),
    .R0_data(mem_253_7_R0_data),
    .R0_en(mem_253_7_R0_en),
    .W0_addr(mem_253_7_W0_addr),
    .W0_clk(mem_253_7_W0_clk),
    .W0_data(mem_253_7_W0_data),
    .W0_en(mem_253_7_W0_en),
    .W0_mask(mem_253_7_W0_mask)
  );
  split_mem_0_ext mem_254_0 (
    .R0_addr(mem_254_0_R0_addr),
    .R0_clk(mem_254_0_R0_clk),
    .R0_data(mem_254_0_R0_data),
    .R0_en(mem_254_0_R0_en),
    .W0_addr(mem_254_0_W0_addr),
    .W0_clk(mem_254_0_W0_clk),
    .W0_data(mem_254_0_W0_data),
    .W0_en(mem_254_0_W0_en),
    .W0_mask(mem_254_0_W0_mask)
  );
  split_mem_0_ext mem_254_1 (
    .R0_addr(mem_254_1_R0_addr),
    .R0_clk(mem_254_1_R0_clk),
    .R0_data(mem_254_1_R0_data),
    .R0_en(mem_254_1_R0_en),
    .W0_addr(mem_254_1_W0_addr),
    .W0_clk(mem_254_1_W0_clk),
    .W0_data(mem_254_1_W0_data),
    .W0_en(mem_254_1_W0_en),
    .W0_mask(mem_254_1_W0_mask)
  );
  split_mem_0_ext mem_254_2 (
    .R0_addr(mem_254_2_R0_addr),
    .R0_clk(mem_254_2_R0_clk),
    .R0_data(mem_254_2_R0_data),
    .R0_en(mem_254_2_R0_en),
    .W0_addr(mem_254_2_W0_addr),
    .W0_clk(mem_254_2_W0_clk),
    .W0_data(mem_254_2_W0_data),
    .W0_en(mem_254_2_W0_en),
    .W0_mask(mem_254_2_W0_mask)
  );
  split_mem_0_ext mem_254_3 (
    .R0_addr(mem_254_3_R0_addr),
    .R0_clk(mem_254_3_R0_clk),
    .R0_data(mem_254_3_R0_data),
    .R0_en(mem_254_3_R0_en),
    .W0_addr(mem_254_3_W0_addr),
    .W0_clk(mem_254_3_W0_clk),
    .W0_data(mem_254_3_W0_data),
    .W0_en(mem_254_3_W0_en),
    .W0_mask(mem_254_3_W0_mask)
  );
  split_mem_0_ext mem_254_4 (
    .R0_addr(mem_254_4_R0_addr),
    .R0_clk(mem_254_4_R0_clk),
    .R0_data(mem_254_4_R0_data),
    .R0_en(mem_254_4_R0_en),
    .W0_addr(mem_254_4_W0_addr),
    .W0_clk(mem_254_4_W0_clk),
    .W0_data(mem_254_4_W0_data),
    .W0_en(mem_254_4_W0_en),
    .W0_mask(mem_254_4_W0_mask)
  );
  split_mem_0_ext mem_254_5 (
    .R0_addr(mem_254_5_R0_addr),
    .R0_clk(mem_254_5_R0_clk),
    .R0_data(mem_254_5_R0_data),
    .R0_en(mem_254_5_R0_en),
    .W0_addr(mem_254_5_W0_addr),
    .W0_clk(mem_254_5_W0_clk),
    .W0_data(mem_254_5_W0_data),
    .W0_en(mem_254_5_W0_en),
    .W0_mask(mem_254_5_W0_mask)
  );
  split_mem_0_ext mem_254_6 (
    .R0_addr(mem_254_6_R0_addr),
    .R0_clk(mem_254_6_R0_clk),
    .R0_data(mem_254_6_R0_data),
    .R0_en(mem_254_6_R0_en),
    .W0_addr(mem_254_6_W0_addr),
    .W0_clk(mem_254_6_W0_clk),
    .W0_data(mem_254_6_W0_data),
    .W0_en(mem_254_6_W0_en),
    .W0_mask(mem_254_6_W0_mask)
  );
  split_mem_0_ext mem_254_7 (
    .R0_addr(mem_254_7_R0_addr),
    .R0_clk(mem_254_7_R0_clk),
    .R0_data(mem_254_7_R0_data),
    .R0_en(mem_254_7_R0_en),
    .W0_addr(mem_254_7_W0_addr),
    .W0_clk(mem_254_7_W0_clk),
    .W0_data(mem_254_7_W0_data),
    .W0_en(mem_254_7_W0_en),
    .W0_mask(mem_254_7_W0_mask)
  );
  split_mem_0_ext mem_255_0 (
    .R0_addr(mem_255_0_R0_addr),
    .R0_clk(mem_255_0_R0_clk),
    .R0_data(mem_255_0_R0_data),
    .R0_en(mem_255_0_R0_en),
    .W0_addr(mem_255_0_W0_addr),
    .W0_clk(mem_255_0_W0_clk),
    .W0_data(mem_255_0_W0_data),
    .W0_en(mem_255_0_W0_en),
    .W0_mask(mem_255_0_W0_mask)
  );
  split_mem_0_ext mem_255_1 (
    .R0_addr(mem_255_1_R0_addr),
    .R0_clk(mem_255_1_R0_clk),
    .R0_data(mem_255_1_R0_data),
    .R0_en(mem_255_1_R0_en),
    .W0_addr(mem_255_1_W0_addr),
    .W0_clk(mem_255_1_W0_clk),
    .W0_data(mem_255_1_W0_data),
    .W0_en(mem_255_1_W0_en),
    .W0_mask(mem_255_1_W0_mask)
  );
  split_mem_0_ext mem_255_2 (
    .R0_addr(mem_255_2_R0_addr),
    .R0_clk(mem_255_2_R0_clk),
    .R0_data(mem_255_2_R0_data),
    .R0_en(mem_255_2_R0_en),
    .W0_addr(mem_255_2_W0_addr),
    .W0_clk(mem_255_2_W0_clk),
    .W0_data(mem_255_2_W0_data),
    .W0_en(mem_255_2_W0_en),
    .W0_mask(mem_255_2_W0_mask)
  );
  split_mem_0_ext mem_255_3 (
    .R0_addr(mem_255_3_R0_addr),
    .R0_clk(mem_255_3_R0_clk),
    .R0_data(mem_255_3_R0_data),
    .R0_en(mem_255_3_R0_en),
    .W0_addr(mem_255_3_W0_addr),
    .W0_clk(mem_255_3_W0_clk),
    .W0_data(mem_255_3_W0_data),
    .W0_en(mem_255_3_W0_en),
    .W0_mask(mem_255_3_W0_mask)
  );
  split_mem_0_ext mem_255_4 (
    .R0_addr(mem_255_4_R0_addr),
    .R0_clk(mem_255_4_R0_clk),
    .R0_data(mem_255_4_R0_data),
    .R0_en(mem_255_4_R0_en),
    .W0_addr(mem_255_4_W0_addr),
    .W0_clk(mem_255_4_W0_clk),
    .W0_data(mem_255_4_W0_data),
    .W0_en(mem_255_4_W0_en),
    .W0_mask(mem_255_4_W0_mask)
  );
  split_mem_0_ext mem_255_5 (
    .R0_addr(mem_255_5_R0_addr),
    .R0_clk(mem_255_5_R0_clk),
    .R0_data(mem_255_5_R0_data),
    .R0_en(mem_255_5_R0_en),
    .W0_addr(mem_255_5_W0_addr),
    .W0_clk(mem_255_5_W0_clk),
    .W0_data(mem_255_5_W0_data),
    .W0_en(mem_255_5_W0_en),
    .W0_mask(mem_255_5_W0_mask)
  );
  split_mem_0_ext mem_255_6 (
    .R0_addr(mem_255_6_R0_addr),
    .R0_clk(mem_255_6_R0_clk),
    .R0_data(mem_255_6_R0_data),
    .R0_en(mem_255_6_R0_en),
    .W0_addr(mem_255_6_W0_addr),
    .W0_clk(mem_255_6_W0_clk),
    .W0_data(mem_255_6_W0_data),
    .W0_en(mem_255_6_W0_en),
    .W0_mask(mem_255_6_W0_mask)
  );
  split_mem_0_ext mem_255_7 (
    .R0_addr(mem_255_7_R0_addr),
    .R0_clk(mem_255_7_R0_clk),
    .R0_data(mem_255_7_R0_data),
    .R0_en(mem_255_7_R0_en),
    .W0_addr(mem_255_7_W0_addr),
    .W0_clk(mem_255_7_W0_clk),
    .W0_data(mem_255_7_W0_data),
    .W0_en(mem_255_7_W0_en),
    .W0_mask(mem_255_7_W0_mask)
  );
  assign R0_data = R0_addr_sel_reg == 8'h0 ? R0_data_0 : R0_addr_sel_reg == 8'h1 ? R0_data_1 : R0_addr_sel_reg == 8'h2
     ? R0_data_2 : R0_addr_sel_reg == 8'h3 ? R0_data_3 : R0_addr_sel_reg == 8'h4 ? R0_data_4 : R0_addr_sel_reg == 8'h5
     ? R0_data_5 : R0_addr_sel_reg == 8'h6 ? R0_data_6 : R0_addr_sel_reg == 8'h7 ? R0_data_7 : R0_addr_sel_reg == 8'h8
     ? R0_data_8 : R0_addr_sel_reg == 8'h9 ? R0_data_9 : R0_addr_sel_reg == 8'ha ? R0_data_10 : R0_addr_sel_reg == 8'hb
     ? R0_data_11 : R0_addr_sel_reg == 8'hc ? R0_data_12 : R0_addr_sel_reg == 8'hd ? R0_data_13 : R0_addr_sel_reg == 8'he
     ? R0_data_14 : R0_addr_sel_reg == 8'hf ? R0_data_15 : R0_addr_sel_reg == 8'h10 ? R0_data_16 : R0_addr_sel_reg == 8'h11
     ? R0_data_17 : R0_addr_sel_reg == 8'h12 ? R0_data_18 : R0_addr_sel_reg == 8'h13 ? R0_data_19 : R0_addr_sel_reg == 8'h14
     ? R0_data_20 : R0_addr_sel_reg == 8'h15 ? R0_data_21 : R0_addr_sel_reg == 8'h16 ? R0_data_22 : R0_addr_sel_reg == 8'h17
     ? R0_data_23 : R0_addr_sel_reg == 8'h18 ? R0_data_24 : R0_addr_sel_reg == 8'h19 ? R0_data_25 : R0_addr_sel_reg == 8'h1a
     ? R0_data_26 : R0_addr_sel_reg == 8'h1b ? R0_data_27 : R0_addr_sel_reg == 8'h1c ? R0_data_28 : R0_addr_sel_reg == 8'h1d
     ? R0_data_29 : R0_addr_sel_reg == 8'h1e ? R0_data_30 : R0_addr_sel_reg == 8'h1f ? R0_data_31 : R0_addr_sel_reg == 8'h20
     ? R0_data_32 : R0_addr_sel_reg == 8'h21 ? R0_data_33 : R0_addr_sel_reg == 8'h22 ? R0_data_34 : R0_addr_sel_reg == 8'h23
     ? R0_data_35 : R0_addr_sel_reg == 8'h24 ? R0_data_36 : R0_addr_sel_reg == 8'h25 ? R0_data_37 : R0_addr_sel_reg == 8'h26
     ? R0_data_38 : R0_addr_sel_reg == 8'h27 ? R0_data_39 : R0_addr_sel_reg == 8'h28 ? R0_data_40 : R0_addr_sel_reg == 8'h29
     ? R0_data_41 : R0_addr_sel_reg == 8'h2a ? R0_data_42 : R0_addr_sel_reg == 8'h2b ? R0_data_43 : R0_addr_sel_reg == 8'h2c
     ? R0_data_44 : R0_addr_sel_reg == 8'h2d ? R0_data_45 : R0_addr_sel_reg == 8'h2e ? R0_data_46 : R0_addr_sel_reg == 8'h2f
     ? R0_data_47 : R0_addr_sel_reg == 8'h30 ? R0_data_48 : R0_addr_sel_reg == 8'h31 ? R0_data_49 : R0_addr_sel_reg == 8'h32
     ? R0_data_50 : R0_addr_sel_reg == 8'h33 ? R0_data_51 : R0_addr_sel_reg == 8'h34 ? R0_data_52 : R0_addr_sel_reg == 8'h35
     ? R0_data_53 : R0_addr_sel_reg == 8'h36 ? R0_data_54 : R0_addr_sel_reg == 8'h37 ? R0_data_55 : R0_addr_sel_reg == 8'h38
     ? R0_data_56 : R0_addr_sel_reg == 8'h39 ? R0_data_57 : R0_addr_sel_reg == 8'h3a ? R0_data_58 : R0_addr_sel_reg == 8'h3b
     ? R0_data_59 : R0_addr_sel_reg == 8'h3c ? R0_data_60 : R0_addr_sel_reg == 8'h3d ? R0_data_61 : R0_addr_sel_reg == 8'h3e
     ? R0_data_62 : R0_addr_sel_reg == 8'h3f ? R0_data_63 : R0_addr_sel_reg == 8'h40 ? R0_data_64 : R0_addr_sel_reg == 8'h41
     ? R0_data_65 : R0_addr_sel_reg == 8'h42 ? R0_data_66 : R0_addr_sel_reg == 8'h43 ? R0_data_67 : R0_addr_sel_reg == 8'h44
     ? R0_data_68 : R0_addr_sel_reg == 8'h45 ? R0_data_69 : R0_addr_sel_reg == 8'h46 ? R0_data_70 : R0_addr_sel_reg == 8'h47
     ? R0_data_71 : R0_addr_sel_reg == 8'h48 ? R0_data_72 : R0_addr_sel_reg == 8'h49 ? R0_data_73 : R0_addr_sel_reg == 8'h4a
     ? R0_data_74 : R0_addr_sel_reg == 8'h4b ? R0_data_75 : R0_addr_sel_reg == 8'h4c ? R0_data_76 : R0_addr_sel_reg == 8'h4d
     ? R0_data_77 : R0_addr_sel_reg == 8'h4e ? R0_data_78 : R0_addr_sel_reg == 8'h4f ? R0_data_79 : R0_addr_sel_reg == 8'h50
     ? R0_data_80 : R0_addr_sel_reg == 8'h51 ? R0_data_81 : R0_addr_sel_reg == 8'h52 ? R0_data_82 : R0_addr_sel_reg == 8'h53
     ? R0_data_83 : R0_addr_sel_reg == 8'h54 ? R0_data_84 : R0_addr_sel_reg == 8'h55 ? R0_data_85 : R0_addr_sel_reg == 8'h56
     ? R0_data_86 : R0_addr_sel_reg == 8'h57 ? R0_data_87 : R0_addr_sel_reg == 8'h58 ? R0_data_88 : R0_addr_sel_reg == 8'h59
     ? R0_data_89 : R0_addr_sel_reg == 8'h5a ? R0_data_90 : R0_addr_sel_reg == 8'h5b ? R0_data_91 : R0_addr_sel_reg == 8'h5c
     ? R0_data_92 : R0_addr_sel_reg == 8'h5d ? R0_data_93 : R0_addr_sel_reg == 8'h5e ? R0_data_94 : R0_addr_sel_reg == 8'h5f
     ? R0_data_95 : R0_addr_sel_reg == 8'h60 ? R0_data_96 : R0_addr_sel_reg == 8'h61 ? R0_data_97 : R0_addr_sel_reg == 8'h62
     ? R0_data_98 : R0_addr_sel_reg == 8'h63 ? R0_data_99 : R0_addr_sel_reg == 8'h64 ? R0_data_100 : R0_addr_sel_reg == 8'h65
     ? R0_data_101 : R0_addr_sel_reg == 8'h66 ? R0_data_102 : R0_addr_sel_reg == 8'h67 ? R0_data_103 : R0_addr_sel_reg
     == 8'h68 ? R0_data_104 : R0_addr_sel_reg == 8'h69 ? R0_data_105 : R0_addr_sel_reg == 8'h6a ? R0_data_106 :
    R0_addr_sel_reg == 8'h6b ? R0_data_107 : R0_addr_sel_reg == 8'h6c ? R0_data_108 : R0_addr_sel_reg == 8'h6d ?
    R0_data_109 : R0_addr_sel_reg == 8'h6e ? R0_data_110 : R0_addr_sel_reg == 8'h6f ? R0_data_111 : R0_addr_sel_reg == 8'h70
     ? R0_data_112 : R0_addr_sel_reg == 8'h71 ? R0_data_113 : R0_addr_sel_reg == 8'h72 ? R0_data_114 : R0_addr_sel_reg
     == 8'h73 ? R0_data_115 : R0_addr_sel_reg == 8'h74 ? R0_data_116 : R0_addr_sel_reg == 8'h75 ? R0_data_117 :
    R0_addr_sel_reg == 8'h76 ? R0_data_118 : R0_addr_sel_reg == 8'h77 ? R0_data_119 : R0_addr_sel_reg == 8'h78 ?
    R0_data_120 : R0_addr_sel_reg == 8'h79 ? R0_data_121 : R0_addr_sel_reg == 8'h7a ? R0_data_122 : R0_addr_sel_reg == 8'h7b
     ? R0_data_123 : R0_addr_sel_reg == 8'h7c ? R0_data_124 : R0_addr_sel_reg == 8'h7d ? R0_data_125 : R0_addr_sel_reg
     == 8'h7e ? R0_data_126 : R0_addr_sel_reg == 8'h7f ? R0_data_127 : R0_addr_sel_reg == 8'h80 ? R0_data_128 :
    R0_addr_sel_reg == 8'h81 ? R0_data_129 : R0_addr_sel_reg == 8'h82 ? R0_data_130 : R0_addr_sel_reg == 8'h83 ?
    R0_data_131 : R0_addr_sel_reg == 8'h84 ? R0_data_132 : R0_addr_sel_reg == 8'h85 ? R0_data_133 : R0_addr_sel_reg == 8'h86
     ? R0_data_134 : R0_addr_sel_reg == 8'h87 ? R0_data_135 : R0_addr_sel_reg == 8'h88 ? R0_data_136 : R0_addr_sel_reg
     == 8'h89 ? R0_data_137 : R0_addr_sel_reg == 8'h8a ? R0_data_138 : R0_addr_sel_reg == 8'h8b ? R0_data_139 :
    R0_addr_sel_reg == 8'h8c ? R0_data_140 : R0_addr_sel_reg == 8'h8d ? R0_data_141 : R0_addr_sel_reg == 8'h8e ?
    R0_data_142 : R0_addr_sel_reg == 8'h8f ? R0_data_143 : R0_addr_sel_reg == 8'h90 ? R0_data_144 : R0_addr_sel_reg == 8'h91
     ? R0_data_145 : R0_addr_sel_reg == 8'h92 ? R0_data_146 : R0_addr_sel_reg == 8'h93 ? R0_data_147 : R0_addr_sel_reg
     == 8'h94 ? R0_data_148 : R0_addr_sel_reg == 8'h95 ? R0_data_149 : R0_addr_sel_reg == 8'h96 ? R0_data_150 :
    R0_addr_sel_reg == 8'h97 ? R0_data_151 : R0_addr_sel_reg == 8'h98 ? R0_data_152 : R0_addr_sel_reg == 8'h99 ?
    R0_data_153 : R0_addr_sel_reg == 8'h9a ? R0_data_154 : R0_addr_sel_reg == 8'h9b ? R0_data_155 : R0_addr_sel_reg == 8'h9c
     ? R0_data_156 : R0_addr_sel_reg == 8'h9d ? R0_data_157 : R0_addr_sel_reg == 8'h9e ? R0_data_158 : R0_addr_sel_reg
     == 8'h9f ? R0_data_159 : R0_addr_sel_reg == 8'ha0 ? R0_data_160 : R0_addr_sel_reg == 8'ha1 ? R0_data_161 :
    R0_addr_sel_reg == 8'ha2 ? R0_data_162 : R0_addr_sel_reg == 8'ha3 ? R0_data_163 : R0_addr_sel_reg == 8'ha4 ?
    R0_data_164 : R0_addr_sel_reg == 8'ha5 ? R0_data_165 : R0_addr_sel_reg == 8'ha6 ? R0_data_166 : R0_addr_sel_reg == 8'ha7
     ? R0_data_167 : R0_addr_sel_reg == 8'ha8 ? R0_data_168 : R0_addr_sel_reg == 8'ha9 ? R0_data_169 : R0_addr_sel_reg
     == 8'haa ? R0_data_170 : R0_addr_sel_reg == 8'hab ? R0_data_171 : R0_addr_sel_reg == 8'hac ? R0_data_172 :
    R0_addr_sel_reg == 8'had ? R0_data_173 : R0_addr_sel_reg == 8'hae ? R0_data_174 : R0_addr_sel_reg == 8'haf ?
    R0_data_175 : R0_addr_sel_reg == 8'hb0 ? R0_data_176 : R0_addr_sel_reg == 8'hb1 ? R0_data_177 : R0_addr_sel_reg == 8'hb2
     ? R0_data_178 : R0_addr_sel_reg == 8'hb3 ? R0_data_179 : R0_addr_sel_reg == 8'hb4 ? R0_data_180 : R0_addr_sel_reg
     == 8'hb5 ? R0_data_181 : R0_addr_sel_reg == 8'hb6 ? R0_data_182 : R0_addr_sel_reg == 8'hb7 ? R0_data_183 :
    R0_addr_sel_reg == 8'hb8 ? R0_data_184 : R0_addr_sel_reg == 8'hb9 ? R0_data_185 : R0_addr_sel_reg == 8'hba ?
    R0_data_186 : R0_addr_sel_reg == 8'hbb ? R0_data_187 : R0_addr_sel_reg == 8'hbc ? R0_data_188 : R0_addr_sel_reg == 8'hbd
     ? R0_data_189 : R0_addr_sel_reg == 8'hbe ? R0_data_190 : R0_addr_sel_reg == 8'hbf ? R0_data_191 : R0_addr_sel_reg
     == 8'hc0 ? R0_data_192 : R0_addr_sel_reg == 8'hc1 ? R0_data_193 : R0_addr_sel_reg == 8'hc2 ? R0_data_194 :
    R0_addr_sel_reg == 8'hc3 ? R0_data_195 : R0_addr_sel_reg == 8'hc4 ? R0_data_196 : R0_addr_sel_reg == 8'hc5 ?
    R0_data_197 : R0_addr_sel_reg == 8'hc6 ? R0_data_198 : R0_addr_sel_reg == 8'hc7 ? R0_data_199 : R0_addr_sel_reg == 8'hc8
     ? R0_data_200 : R0_addr_sel_reg == 8'hc9 ? R0_data_201 : R0_addr_sel_reg == 8'hca ? R0_data_202 : R0_addr_sel_reg
     == 8'hcb ? R0_data_203 : R0_addr_sel_reg == 8'hcc ? R0_data_204 : R0_addr_sel_reg == 8'hcd ? R0_data_205 :
    R0_addr_sel_reg == 8'hce ? R0_data_206 : R0_addr_sel_reg == 8'hcf ? R0_data_207 : R0_addr_sel_reg == 8'hd0 ?
    R0_data_208 : R0_addr_sel_reg == 8'hd1 ? R0_data_209 : R0_addr_sel_reg == 8'hd2 ? R0_data_210 : R0_addr_sel_reg == 8'hd3
     ? R0_data_211 : R0_addr_sel_reg == 8'hd4 ? R0_data_212 : R0_addr_sel_reg == 8'hd5 ? R0_data_213 : R0_addr_sel_reg
     == 8'hd6 ? R0_data_214 : R0_addr_sel_reg == 8'hd7 ? R0_data_215 : R0_addr_sel_reg == 8'hd8 ? R0_data_216 :
    R0_addr_sel_reg == 8'hd9 ? R0_data_217 : R0_addr_sel_reg == 8'hda ? R0_data_218 : R0_addr_sel_reg == 8'hdb ?
    R0_data_219 : R0_addr_sel_reg == 8'hdc ? R0_data_220 : R0_addr_sel_reg == 8'hdd ? R0_data_221 : R0_addr_sel_reg == 8'hde
     ? R0_data_222 : R0_addr_sel_reg == 8'hdf ? R0_data_223 : R0_addr_sel_reg == 8'he0 ? R0_data_224 : R0_addr_sel_reg
     == 8'he1 ? R0_data_225 : R0_addr_sel_reg == 8'he2 ? R0_data_226 : R0_addr_sel_reg == 8'he3 ? R0_data_227 :
    R0_addr_sel_reg == 8'he4 ? R0_data_228 : R0_addr_sel_reg == 8'he5 ? R0_data_229 : R0_addr_sel_reg == 8'he6 ?
    R0_data_230 : R0_addr_sel_reg == 8'he7 ? R0_data_231 : R0_addr_sel_reg == 8'he8 ? R0_data_232 : R0_addr_sel_reg == 8'he9
     ? R0_data_233 : R0_addr_sel_reg == 8'hea ? R0_data_234 : R0_addr_sel_reg == 8'heb ? R0_data_235 : R0_addr_sel_reg
     == 8'hec ? R0_data_236 : R0_addr_sel_reg == 8'hed ? R0_data_237 : R0_addr_sel_reg == 8'hee ? R0_data_238 :
    R0_addr_sel_reg == 8'hef ? R0_data_239 : R0_addr_sel_reg == 8'hf0 ? R0_data_240 : R0_addr_sel_reg == 8'hf1 ?
    R0_data_241 : R0_addr_sel_reg == 8'hf2 ? R0_data_242 : R0_addr_sel_reg == 8'hf3 ? R0_data_243 : R0_addr_sel_reg == 8'hf4
     ? R0_data_244 : R0_addr_sel_reg == 8'hf5 ? R0_data_245 : R0_addr_sel_reg == 8'hf6 ? R0_data_246 : R0_addr_sel_reg
     == 8'hf7 ? R0_data_247 : R0_addr_sel_reg == 8'hf8 ? R0_data_248 : R0_addr_sel_reg == 8'hf9 ? R0_data_249 :
    R0_addr_sel_reg == 8'hfa ? R0_data_250 : R0_addr_sel_reg == 8'hfb ? R0_data_251 : R0_addr_sel_reg == 8'hfc ?
    R0_data_252 : R0_addr_sel_reg == 8'hfd ? R0_data_253 : R0_addr_sel_reg == 8'hfe ? R0_data_254 : R0_addr_sel_reg == 8'hff
     ? R0_data_255 : 64'h0;
  assign mem_0_0_R0_addr = R0_addr[25:0];
  assign mem_0_0_R0_clk = R0_clk;
  assign mem_0_0_R0_en = R0_en & R0_addr_sel == 8'h0;
  assign mem_0_0_W0_addr = W0_addr[25:0];
  assign mem_0_0_W0_clk = W0_clk;
  assign mem_0_0_W0_data = W0_data[7:0];
  assign mem_0_0_W0_en = W0_en & W0_addr_sel == 8'h0;
  assign mem_0_0_W0_mask = W0_mask[0];
  assign mem_0_1_R0_addr = R0_addr[25:0];
  assign mem_0_1_R0_clk = R0_clk;
  assign mem_0_1_R0_en = R0_en & R0_addr_sel == 8'h0;
  assign mem_0_1_W0_addr = W0_addr[25:0];
  assign mem_0_1_W0_clk = W0_clk;
  assign mem_0_1_W0_data = W0_data[15:8];
  assign mem_0_1_W0_en = W0_en & W0_addr_sel == 8'h0;
  assign mem_0_1_W0_mask = W0_mask[1];
  assign mem_0_2_R0_addr = R0_addr[25:0];
  assign mem_0_2_R0_clk = R0_clk;
  assign mem_0_2_R0_en = R0_en & R0_addr_sel == 8'h0;
  assign mem_0_2_W0_addr = W0_addr[25:0];
  assign mem_0_2_W0_clk = W0_clk;
  assign mem_0_2_W0_data = W0_data[23:16];
  assign mem_0_2_W0_en = W0_en & W0_addr_sel == 8'h0;
  assign mem_0_2_W0_mask = W0_mask[2];
  assign mem_0_3_R0_addr = R0_addr[25:0];
  assign mem_0_3_R0_clk = R0_clk;
  assign mem_0_3_R0_en = R0_en & R0_addr_sel == 8'h0;
  assign mem_0_3_W0_addr = W0_addr[25:0];
  assign mem_0_3_W0_clk = W0_clk;
  assign mem_0_3_W0_data = W0_data[31:24];
  assign mem_0_3_W0_en = W0_en & W0_addr_sel == 8'h0;
  assign mem_0_3_W0_mask = W0_mask[3];
  assign mem_0_4_R0_addr = R0_addr[25:0];
  assign mem_0_4_R0_clk = R0_clk;
  assign mem_0_4_R0_en = R0_en & R0_addr_sel == 8'h0;
  assign mem_0_4_W0_addr = W0_addr[25:0];
  assign mem_0_4_W0_clk = W0_clk;
  assign mem_0_4_W0_data = W0_data[39:32];
  assign mem_0_4_W0_en = W0_en & W0_addr_sel == 8'h0;
  assign mem_0_4_W0_mask = W0_mask[4];
  assign mem_0_5_R0_addr = R0_addr[25:0];
  assign mem_0_5_R0_clk = R0_clk;
  assign mem_0_5_R0_en = R0_en & R0_addr_sel == 8'h0;
  assign mem_0_5_W0_addr = W0_addr[25:0];
  assign mem_0_5_W0_clk = W0_clk;
  assign mem_0_5_W0_data = W0_data[47:40];
  assign mem_0_5_W0_en = W0_en & W0_addr_sel == 8'h0;
  assign mem_0_5_W0_mask = W0_mask[5];
  assign mem_0_6_R0_addr = R0_addr[25:0];
  assign mem_0_6_R0_clk = R0_clk;
  assign mem_0_6_R0_en = R0_en & R0_addr_sel == 8'h0;
  assign mem_0_6_W0_addr = W0_addr[25:0];
  assign mem_0_6_W0_clk = W0_clk;
  assign mem_0_6_W0_data = W0_data[55:48];
  assign mem_0_6_W0_en = W0_en & W0_addr_sel == 8'h0;
  assign mem_0_6_W0_mask = W0_mask[6];
  assign mem_0_7_R0_addr = R0_addr[25:0];
  assign mem_0_7_R0_clk = R0_clk;
  assign mem_0_7_R0_en = R0_en & R0_addr_sel == 8'h0;
  assign mem_0_7_W0_addr = W0_addr[25:0];
  assign mem_0_7_W0_clk = W0_clk;
  assign mem_0_7_W0_data = W0_data[63:56];
  assign mem_0_7_W0_en = W0_en & W0_addr_sel == 8'h0;
  assign mem_0_7_W0_mask = W0_mask[7];
  assign mem_1_0_R0_addr = R0_addr[25:0];
  assign mem_1_0_R0_clk = R0_clk;
  assign mem_1_0_R0_en = R0_en & R0_addr_sel == 8'h1;
  assign mem_1_0_W0_addr = W0_addr[25:0];
  assign mem_1_0_W0_clk = W0_clk;
  assign mem_1_0_W0_data = W0_data[7:0];
  assign mem_1_0_W0_en = W0_en & W0_addr_sel == 8'h1;
  assign mem_1_0_W0_mask = W0_mask[0];
  assign mem_1_1_R0_addr = R0_addr[25:0];
  assign mem_1_1_R0_clk = R0_clk;
  assign mem_1_1_R0_en = R0_en & R0_addr_sel == 8'h1;
  assign mem_1_1_W0_addr = W0_addr[25:0];
  assign mem_1_1_W0_clk = W0_clk;
  assign mem_1_1_W0_data = W0_data[15:8];
  assign mem_1_1_W0_en = W0_en & W0_addr_sel == 8'h1;
  assign mem_1_1_W0_mask = W0_mask[1];
  assign mem_1_2_R0_addr = R0_addr[25:0];
  assign mem_1_2_R0_clk = R0_clk;
  assign mem_1_2_R0_en = R0_en & R0_addr_sel == 8'h1;
  assign mem_1_2_W0_addr = W0_addr[25:0];
  assign mem_1_2_W0_clk = W0_clk;
  assign mem_1_2_W0_data = W0_data[23:16];
  assign mem_1_2_W0_en = W0_en & W0_addr_sel == 8'h1;
  assign mem_1_2_W0_mask = W0_mask[2];
  assign mem_1_3_R0_addr = R0_addr[25:0];
  assign mem_1_3_R0_clk = R0_clk;
  assign mem_1_3_R0_en = R0_en & R0_addr_sel == 8'h1;
  assign mem_1_3_W0_addr = W0_addr[25:0];
  assign mem_1_3_W0_clk = W0_clk;
  assign mem_1_3_W0_data = W0_data[31:24];
  assign mem_1_3_W0_en = W0_en & W0_addr_sel == 8'h1;
  assign mem_1_3_W0_mask = W0_mask[3];
  assign mem_1_4_R0_addr = R0_addr[25:0];
  assign mem_1_4_R0_clk = R0_clk;
  assign mem_1_4_R0_en = R0_en & R0_addr_sel == 8'h1;
  assign mem_1_4_W0_addr = W0_addr[25:0];
  assign mem_1_4_W0_clk = W0_clk;
  assign mem_1_4_W0_data = W0_data[39:32];
  assign mem_1_4_W0_en = W0_en & W0_addr_sel == 8'h1;
  assign mem_1_4_W0_mask = W0_mask[4];
  assign mem_1_5_R0_addr = R0_addr[25:0];
  assign mem_1_5_R0_clk = R0_clk;
  assign mem_1_5_R0_en = R0_en & R0_addr_sel == 8'h1;
  assign mem_1_5_W0_addr = W0_addr[25:0];
  assign mem_1_5_W0_clk = W0_clk;
  assign mem_1_5_W0_data = W0_data[47:40];
  assign mem_1_5_W0_en = W0_en & W0_addr_sel == 8'h1;
  assign mem_1_5_W0_mask = W0_mask[5];
  assign mem_1_6_R0_addr = R0_addr[25:0];
  assign mem_1_6_R0_clk = R0_clk;
  assign mem_1_6_R0_en = R0_en & R0_addr_sel == 8'h1;
  assign mem_1_6_W0_addr = W0_addr[25:0];
  assign mem_1_6_W0_clk = W0_clk;
  assign mem_1_6_W0_data = W0_data[55:48];
  assign mem_1_6_W0_en = W0_en & W0_addr_sel == 8'h1;
  assign mem_1_6_W0_mask = W0_mask[6];
  assign mem_1_7_R0_addr = R0_addr[25:0];
  assign mem_1_7_R0_clk = R0_clk;
  assign mem_1_7_R0_en = R0_en & R0_addr_sel == 8'h1;
  assign mem_1_7_W0_addr = W0_addr[25:0];
  assign mem_1_7_W0_clk = W0_clk;
  assign mem_1_7_W0_data = W0_data[63:56];
  assign mem_1_7_W0_en = W0_en & W0_addr_sel == 8'h1;
  assign mem_1_7_W0_mask = W0_mask[7];
  assign mem_2_0_R0_addr = R0_addr[25:0];
  assign mem_2_0_R0_clk = R0_clk;
  assign mem_2_0_R0_en = R0_en & R0_addr_sel == 8'h2;
  assign mem_2_0_W0_addr = W0_addr[25:0];
  assign mem_2_0_W0_clk = W0_clk;
  assign mem_2_0_W0_data = W0_data[7:0];
  assign mem_2_0_W0_en = W0_en & W0_addr_sel == 8'h2;
  assign mem_2_0_W0_mask = W0_mask[0];
  assign mem_2_1_R0_addr = R0_addr[25:0];
  assign mem_2_1_R0_clk = R0_clk;
  assign mem_2_1_R0_en = R0_en & R0_addr_sel == 8'h2;
  assign mem_2_1_W0_addr = W0_addr[25:0];
  assign mem_2_1_W0_clk = W0_clk;
  assign mem_2_1_W0_data = W0_data[15:8];
  assign mem_2_1_W0_en = W0_en & W0_addr_sel == 8'h2;
  assign mem_2_1_W0_mask = W0_mask[1];
  assign mem_2_2_R0_addr = R0_addr[25:0];
  assign mem_2_2_R0_clk = R0_clk;
  assign mem_2_2_R0_en = R0_en & R0_addr_sel == 8'h2;
  assign mem_2_2_W0_addr = W0_addr[25:0];
  assign mem_2_2_W0_clk = W0_clk;
  assign mem_2_2_W0_data = W0_data[23:16];
  assign mem_2_2_W0_en = W0_en & W0_addr_sel == 8'h2;
  assign mem_2_2_W0_mask = W0_mask[2];
  assign mem_2_3_R0_addr = R0_addr[25:0];
  assign mem_2_3_R0_clk = R0_clk;
  assign mem_2_3_R0_en = R0_en & R0_addr_sel == 8'h2;
  assign mem_2_3_W0_addr = W0_addr[25:0];
  assign mem_2_3_W0_clk = W0_clk;
  assign mem_2_3_W0_data = W0_data[31:24];
  assign mem_2_3_W0_en = W0_en & W0_addr_sel == 8'h2;
  assign mem_2_3_W0_mask = W0_mask[3];
  assign mem_2_4_R0_addr = R0_addr[25:0];
  assign mem_2_4_R0_clk = R0_clk;
  assign mem_2_4_R0_en = R0_en & R0_addr_sel == 8'h2;
  assign mem_2_4_W0_addr = W0_addr[25:0];
  assign mem_2_4_W0_clk = W0_clk;
  assign mem_2_4_W0_data = W0_data[39:32];
  assign mem_2_4_W0_en = W0_en & W0_addr_sel == 8'h2;
  assign mem_2_4_W0_mask = W0_mask[4];
  assign mem_2_5_R0_addr = R0_addr[25:0];
  assign mem_2_5_R0_clk = R0_clk;
  assign mem_2_5_R0_en = R0_en & R0_addr_sel == 8'h2;
  assign mem_2_5_W0_addr = W0_addr[25:0];
  assign mem_2_5_W0_clk = W0_clk;
  assign mem_2_5_W0_data = W0_data[47:40];
  assign mem_2_5_W0_en = W0_en & W0_addr_sel == 8'h2;
  assign mem_2_5_W0_mask = W0_mask[5];
  assign mem_2_6_R0_addr = R0_addr[25:0];
  assign mem_2_6_R0_clk = R0_clk;
  assign mem_2_6_R0_en = R0_en & R0_addr_sel == 8'h2;
  assign mem_2_6_W0_addr = W0_addr[25:0];
  assign mem_2_6_W0_clk = W0_clk;
  assign mem_2_6_W0_data = W0_data[55:48];
  assign mem_2_6_W0_en = W0_en & W0_addr_sel == 8'h2;
  assign mem_2_6_W0_mask = W0_mask[6];
  assign mem_2_7_R0_addr = R0_addr[25:0];
  assign mem_2_7_R0_clk = R0_clk;
  assign mem_2_7_R0_en = R0_en & R0_addr_sel == 8'h2;
  assign mem_2_7_W0_addr = W0_addr[25:0];
  assign mem_2_7_W0_clk = W0_clk;
  assign mem_2_7_W0_data = W0_data[63:56];
  assign mem_2_7_W0_en = W0_en & W0_addr_sel == 8'h2;
  assign mem_2_7_W0_mask = W0_mask[7];
  assign mem_3_0_R0_addr = R0_addr[25:0];
  assign mem_3_0_R0_clk = R0_clk;
  assign mem_3_0_R0_en = R0_en & R0_addr_sel == 8'h3;
  assign mem_3_0_W0_addr = W0_addr[25:0];
  assign mem_3_0_W0_clk = W0_clk;
  assign mem_3_0_W0_data = W0_data[7:0];
  assign mem_3_0_W0_en = W0_en & W0_addr_sel == 8'h3;
  assign mem_3_0_W0_mask = W0_mask[0];
  assign mem_3_1_R0_addr = R0_addr[25:0];
  assign mem_3_1_R0_clk = R0_clk;
  assign mem_3_1_R0_en = R0_en & R0_addr_sel == 8'h3;
  assign mem_3_1_W0_addr = W0_addr[25:0];
  assign mem_3_1_W0_clk = W0_clk;
  assign mem_3_1_W0_data = W0_data[15:8];
  assign mem_3_1_W0_en = W0_en & W0_addr_sel == 8'h3;
  assign mem_3_1_W0_mask = W0_mask[1];
  assign mem_3_2_R0_addr = R0_addr[25:0];
  assign mem_3_2_R0_clk = R0_clk;
  assign mem_3_2_R0_en = R0_en & R0_addr_sel == 8'h3;
  assign mem_3_2_W0_addr = W0_addr[25:0];
  assign mem_3_2_W0_clk = W0_clk;
  assign mem_3_2_W0_data = W0_data[23:16];
  assign mem_3_2_W0_en = W0_en & W0_addr_sel == 8'h3;
  assign mem_3_2_W0_mask = W0_mask[2];
  assign mem_3_3_R0_addr = R0_addr[25:0];
  assign mem_3_3_R0_clk = R0_clk;
  assign mem_3_3_R0_en = R0_en & R0_addr_sel == 8'h3;
  assign mem_3_3_W0_addr = W0_addr[25:0];
  assign mem_3_3_W0_clk = W0_clk;
  assign mem_3_3_W0_data = W0_data[31:24];
  assign mem_3_3_W0_en = W0_en & W0_addr_sel == 8'h3;
  assign mem_3_3_W0_mask = W0_mask[3];
  assign mem_3_4_R0_addr = R0_addr[25:0];
  assign mem_3_4_R0_clk = R0_clk;
  assign mem_3_4_R0_en = R0_en & R0_addr_sel == 8'h3;
  assign mem_3_4_W0_addr = W0_addr[25:0];
  assign mem_3_4_W0_clk = W0_clk;
  assign mem_3_4_W0_data = W0_data[39:32];
  assign mem_3_4_W0_en = W0_en & W0_addr_sel == 8'h3;
  assign mem_3_4_W0_mask = W0_mask[4];
  assign mem_3_5_R0_addr = R0_addr[25:0];
  assign mem_3_5_R0_clk = R0_clk;
  assign mem_3_5_R0_en = R0_en & R0_addr_sel == 8'h3;
  assign mem_3_5_W0_addr = W0_addr[25:0];
  assign mem_3_5_W0_clk = W0_clk;
  assign mem_3_5_W0_data = W0_data[47:40];
  assign mem_3_5_W0_en = W0_en & W0_addr_sel == 8'h3;
  assign mem_3_5_W0_mask = W0_mask[5];
  assign mem_3_6_R0_addr = R0_addr[25:0];
  assign mem_3_6_R0_clk = R0_clk;
  assign mem_3_6_R0_en = R0_en & R0_addr_sel == 8'h3;
  assign mem_3_6_W0_addr = W0_addr[25:0];
  assign mem_3_6_W0_clk = W0_clk;
  assign mem_3_6_W0_data = W0_data[55:48];
  assign mem_3_6_W0_en = W0_en & W0_addr_sel == 8'h3;
  assign mem_3_6_W0_mask = W0_mask[6];
  assign mem_3_7_R0_addr = R0_addr[25:0];
  assign mem_3_7_R0_clk = R0_clk;
  assign mem_3_7_R0_en = R0_en & R0_addr_sel == 8'h3;
  assign mem_3_7_W0_addr = W0_addr[25:0];
  assign mem_3_7_W0_clk = W0_clk;
  assign mem_3_7_W0_data = W0_data[63:56];
  assign mem_3_7_W0_en = W0_en & W0_addr_sel == 8'h3;
  assign mem_3_7_W0_mask = W0_mask[7];
  assign mem_4_0_R0_addr = R0_addr[25:0];
  assign mem_4_0_R0_clk = R0_clk;
  assign mem_4_0_R0_en = R0_en & R0_addr_sel == 8'h4;
  assign mem_4_0_W0_addr = W0_addr[25:0];
  assign mem_4_0_W0_clk = W0_clk;
  assign mem_4_0_W0_data = W0_data[7:0];
  assign mem_4_0_W0_en = W0_en & W0_addr_sel == 8'h4;
  assign mem_4_0_W0_mask = W0_mask[0];
  assign mem_4_1_R0_addr = R0_addr[25:0];
  assign mem_4_1_R0_clk = R0_clk;
  assign mem_4_1_R0_en = R0_en & R0_addr_sel == 8'h4;
  assign mem_4_1_W0_addr = W0_addr[25:0];
  assign mem_4_1_W0_clk = W0_clk;
  assign mem_4_1_W0_data = W0_data[15:8];
  assign mem_4_1_W0_en = W0_en & W0_addr_sel == 8'h4;
  assign mem_4_1_W0_mask = W0_mask[1];
  assign mem_4_2_R0_addr = R0_addr[25:0];
  assign mem_4_2_R0_clk = R0_clk;
  assign mem_4_2_R0_en = R0_en & R0_addr_sel == 8'h4;
  assign mem_4_2_W0_addr = W0_addr[25:0];
  assign mem_4_2_W0_clk = W0_clk;
  assign mem_4_2_W0_data = W0_data[23:16];
  assign mem_4_2_W0_en = W0_en & W0_addr_sel == 8'h4;
  assign mem_4_2_W0_mask = W0_mask[2];
  assign mem_4_3_R0_addr = R0_addr[25:0];
  assign mem_4_3_R0_clk = R0_clk;
  assign mem_4_3_R0_en = R0_en & R0_addr_sel == 8'h4;
  assign mem_4_3_W0_addr = W0_addr[25:0];
  assign mem_4_3_W0_clk = W0_clk;
  assign mem_4_3_W0_data = W0_data[31:24];
  assign mem_4_3_W0_en = W0_en & W0_addr_sel == 8'h4;
  assign mem_4_3_W0_mask = W0_mask[3];
  assign mem_4_4_R0_addr = R0_addr[25:0];
  assign mem_4_4_R0_clk = R0_clk;
  assign mem_4_4_R0_en = R0_en & R0_addr_sel == 8'h4;
  assign mem_4_4_W0_addr = W0_addr[25:0];
  assign mem_4_4_W0_clk = W0_clk;
  assign mem_4_4_W0_data = W0_data[39:32];
  assign mem_4_4_W0_en = W0_en & W0_addr_sel == 8'h4;
  assign mem_4_4_W0_mask = W0_mask[4];
  assign mem_4_5_R0_addr = R0_addr[25:0];
  assign mem_4_5_R0_clk = R0_clk;
  assign mem_4_5_R0_en = R0_en & R0_addr_sel == 8'h4;
  assign mem_4_5_W0_addr = W0_addr[25:0];
  assign mem_4_5_W0_clk = W0_clk;
  assign mem_4_5_W0_data = W0_data[47:40];
  assign mem_4_5_W0_en = W0_en & W0_addr_sel == 8'h4;
  assign mem_4_5_W0_mask = W0_mask[5];
  assign mem_4_6_R0_addr = R0_addr[25:0];
  assign mem_4_6_R0_clk = R0_clk;
  assign mem_4_6_R0_en = R0_en & R0_addr_sel == 8'h4;
  assign mem_4_6_W0_addr = W0_addr[25:0];
  assign mem_4_6_W0_clk = W0_clk;
  assign mem_4_6_W0_data = W0_data[55:48];
  assign mem_4_6_W0_en = W0_en & W0_addr_sel == 8'h4;
  assign mem_4_6_W0_mask = W0_mask[6];
  assign mem_4_7_R0_addr = R0_addr[25:0];
  assign mem_4_7_R0_clk = R0_clk;
  assign mem_4_7_R0_en = R0_en & R0_addr_sel == 8'h4;
  assign mem_4_7_W0_addr = W0_addr[25:0];
  assign mem_4_7_W0_clk = W0_clk;
  assign mem_4_7_W0_data = W0_data[63:56];
  assign mem_4_7_W0_en = W0_en & W0_addr_sel == 8'h4;
  assign mem_4_7_W0_mask = W0_mask[7];
  assign mem_5_0_R0_addr = R0_addr[25:0];
  assign mem_5_0_R0_clk = R0_clk;
  assign mem_5_0_R0_en = R0_en & R0_addr_sel == 8'h5;
  assign mem_5_0_W0_addr = W0_addr[25:0];
  assign mem_5_0_W0_clk = W0_clk;
  assign mem_5_0_W0_data = W0_data[7:0];
  assign mem_5_0_W0_en = W0_en & W0_addr_sel == 8'h5;
  assign mem_5_0_W0_mask = W0_mask[0];
  assign mem_5_1_R0_addr = R0_addr[25:0];
  assign mem_5_1_R0_clk = R0_clk;
  assign mem_5_1_R0_en = R0_en & R0_addr_sel == 8'h5;
  assign mem_5_1_W0_addr = W0_addr[25:0];
  assign mem_5_1_W0_clk = W0_clk;
  assign mem_5_1_W0_data = W0_data[15:8];
  assign mem_5_1_W0_en = W0_en & W0_addr_sel == 8'h5;
  assign mem_5_1_W0_mask = W0_mask[1];
  assign mem_5_2_R0_addr = R0_addr[25:0];
  assign mem_5_2_R0_clk = R0_clk;
  assign mem_5_2_R0_en = R0_en & R0_addr_sel == 8'h5;
  assign mem_5_2_W0_addr = W0_addr[25:0];
  assign mem_5_2_W0_clk = W0_clk;
  assign mem_5_2_W0_data = W0_data[23:16];
  assign mem_5_2_W0_en = W0_en & W0_addr_sel == 8'h5;
  assign mem_5_2_W0_mask = W0_mask[2];
  assign mem_5_3_R0_addr = R0_addr[25:0];
  assign mem_5_3_R0_clk = R0_clk;
  assign mem_5_3_R0_en = R0_en & R0_addr_sel == 8'h5;
  assign mem_5_3_W0_addr = W0_addr[25:0];
  assign mem_5_3_W0_clk = W0_clk;
  assign mem_5_3_W0_data = W0_data[31:24];
  assign mem_5_3_W0_en = W0_en & W0_addr_sel == 8'h5;
  assign mem_5_3_W0_mask = W0_mask[3];
  assign mem_5_4_R0_addr = R0_addr[25:0];
  assign mem_5_4_R0_clk = R0_clk;
  assign mem_5_4_R0_en = R0_en & R0_addr_sel == 8'h5;
  assign mem_5_4_W0_addr = W0_addr[25:0];
  assign mem_5_4_W0_clk = W0_clk;
  assign mem_5_4_W0_data = W0_data[39:32];
  assign mem_5_4_W0_en = W0_en & W0_addr_sel == 8'h5;
  assign mem_5_4_W0_mask = W0_mask[4];
  assign mem_5_5_R0_addr = R0_addr[25:0];
  assign mem_5_5_R0_clk = R0_clk;
  assign mem_5_5_R0_en = R0_en & R0_addr_sel == 8'h5;
  assign mem_5_5_W0_addr = W0_addr[25:0];
  assign mem_5_5_W0_clk = W0_clk;
  assign mem_5_5_W0_data = W0_data[47:40];
  assign mem_5_5_W0_en = W0_en & W0_addr_sel == 8'h5;
  assign mem_5_5_W0_mask = W0_mask[5];
  assign mem_5_6_R0_addr = R0_addr[25:0];
  assign mem_5_6_R0_clk = R0_clk;
  assign mem_5_6_R0_en = R0_en & R0_addr_sel == 8'h5;
  assign mem_5_6_W0_addr = W0_addr[25:0];
  assign mem_5_6_W0_clk = W0_clk;
  assign mem_5_6_W0_data = W0_data[55:48];
  assign mem_5_6_W0_en = W0_en & W0_addr_sel == 8'h5;
  assign mem_5_6_W0_mask = W0_mask[6];
  assign mem_5_7_R0_addr = R0_addr[25:0];
  assign mem_5_7_R0_clk = R0_clk;
  assign mem_5_7_R0_en = R0_en & R0_addr_sel == 8'h5;
  assign mem_5_7_W0_addr = W0_addr[25:0];
  assign mem_5_7_W0_clk = W0_clk;
  assign mem_5_7_W0_data = W0_data[63:56];
  assign mem_5_7_W0_en = W0_en & W0_addr_sel == 8'h5;
  assign mem_5_7_W0_mask = W0_mask[7];
  assign mem_6_0_R0_addr = R0_addr[25:0];
  assign mem_6_0_R0_clk = R0_clk;
  assign mem_6_0_R0_en = R0_en & R0_addr_sel == 8'h6;
  assign mem_6_0_W0_addr = W0_addr[25:0];
  assign mem_6_0_W0_clk = W0_clk;
  assign mem_6_0_W0_data = W0_data[7:0];
  assign mem_6_0_W0_en = W0_en & W0_addr_sel == 8'h6;
  assign mem_6_0_W0_mask = W0_mask[0];
  assign mem_6_1_R0_addr = R0_addr[25:0];
  assign mem_6_1_R0_clk = R0_clk;
  assign mem_6_1_R0_en = R0_en & R0_addr_sel == 8'h6;
  assign mem_6_1_W0_addr = W0_addr[25:0];
  assign mem_6_1_W0_clk = W0_clk;
  assign mem_6_1_W0_data = W0_data[15:8];
  assign mem_6_1_W0_en = W0_en & W0_addr_sel == 8'h6;
  assign mem_6_1_W0_mask = W0_mask[1];
  assign mem_6_2_R0_addr = R0_addr[25:0];
  assign mem_6_2_R0_clk = R0_clk;
  assign mem_6_2_R0_en = R0_en & R0_addr_sel == 8'h6;
  assign mem_6_2_W0_addr = W0_addr[25:0];
  assign mem_6_2_W0_clk = W0_clk;
  assign mem_6_2_W0_data = W0_data[23:16];
  assign mem_6_2_W0_en = W0_en & W0_addr_sel == 8'h6;
  assign mem_6_2_W0_mask = W0_mask[2];
  assign mem_6_3_R0_addr = R0_addr[25:0];
  assign mem_6_3_R0_clk = R0_clk;
  assign mem_6_3_R0_en = R0_en & R0_addr_sel == 8'h6;
  assign mem_6_3_W0_addr = W0_addr[25:0];
  assign mem_6_3_W0_clk = W0_clk;
  assign mem_6_3_W0_data = W0_data[31:24];
  assign mem_6_3_W0_en = W0_en & W0_addr_sel == 8'h6;
  assign mem_6_3_W0_mask = W0_mask[3];
  assign mem_6_4_R0_addr = R0_addr[25:0];
  assign mem_6_4_R0_clk = R0_clk;
  assign mem_6_4_R0_en = R0_en & R0_addr_sel == 8'h6;
  assign mem_6_4_W0_addr = W0_addr[25:0];
  assign mem_6_4_W0_clk = W0_clk;
  assign mem_6_4_W0_data = W0_data[39:32];
  assign mem_6_4_W0_en = W0_en & W0_addr_sel == 8'h6;
  assign mem_6_4_W0_mask = W0_mask[4];
  assign mem_6_5_R0_addr = R0_addr[25:0];
  assign mem_6_5_R0_clk = R0_clk;
  assign mem_6_5_R0_en = R0_en & R0_addr_sel == 8'h6;
  assign mem_6_5_W0_addr = W0_addr[25:0];
  assign mem_6_5_W0_clk = W0_clk;
  assign mem_6_5_W0_data = W0_data[47:40];
  assign mem_6_5_W0_en = W0_en & W0_addr_sel == 8'h6;
  assign mem_6_5_W0_mask = W0_mask[5];
  assign mem_6_6_R0_addr = R0_addr[25:0];
  assign mem_6_6_R0_clk = R0_clk;
  assign mem_6_6_R0_en = R0_en & R0_addr_sel == 8'h6;
  assign mem_6_6_W0_addr = W0_addr[25:0];
  assign mem_6_6_W0_clk = W0_clk;
  assign mem_6_6_W0_data = W0_data[55:48];
  assign mem_6_6_W0_en = W0_en & W0_addr_sel == 8'h6;
  assign mem_6_6_W0_mask = W0_mask[6];
  assign mem_6_7_R0_addr = R0_addr[25:0];
  assign mem_6_7_R0_clk = R0_clk;
  assign mem_6_7_R0_en = R0_en & R0_addr_sel == 8'h6;
  assign mem_6_7_W0_addr = W0_addr[25:0];
  assign mem_6_7_W0_clk = W0_clk;
  assign mem_6_7_W0_data = W0_data[63:56];
  assign mem_6_7_W0_en = W0_en & W0_addr_sel == 8'h6;
  assign mem_6_7_W0_mask = W0_mask[7];
  assign mem_7_0_R0_addr = R0_addr[25:0];
  assign mem_7_0_R0_clk = R0_clk;
  assign mem_7_0_R0_en = R0_en & R0_addr_sel == 8'h7;
  assign mem_7_0_W0_addr = W0_addr[25:0];
  assign mem_7_0_W0_clk = W0_clk;
  assign mem_7_0_W0_data = W0_data[7:0];
  assign mem_7_0_W0_en = W0_en & W0_addr_sel == 8'h7;
  assign mem_7_0_W0_mask = W0_mask[0];
  assign mem_7_1_R0_addr = R0_addr[25:0];
  assign mem_7_1_R0_clk = R0_clk;
  assign mem_7_1_R0_en = R0_en & R0_addr_sel == 8'h7;
  assign mem_7_1_W0_addr = W0_addr[25:0];
  assign mem_7_1_W0_clk = W0_clk;
  assign mem_7_1_W0_data = W0_data[15:8];
  assign mem_7_1_W0_en = W0_en & W0_addr_sel == 8'h7;
  assign mem_7_1_W0_mask = W0_mask[1];
  assign mem_7_2_R0_addr = R0_addr[25:0];
  assign mem_7_2_R0_clk = R0_clk;
  assign mem_7_2_R0_en = R0_en & R0_addr_sel == 8'h7;
  assign mem_7_2_W0_addr = W0_addr[25:0];
  assign mem_7_2_W0_clk = W0_clk;
  assign mem_7_2_W0_data = W0_data[23:16];
  assign mem_7_2_W0_en = W0_en & W0_addr_sel == 8'h7;
  assign mem_7_2_W0_mask = W0_mask[2];
  assign mem_7_3_R0_addr = R0_addr[25:0];
  assign mem_7_3_R0_clk = R0_clk;
  assign mem_7_3_R0_en = R0_en & R0_addr_sel == 8'h7;
  assign mem_7_3_W0_addr = W0_addr[25:0];
  assign mem_7_3_W0_clk = W0_clk;
  assign mem_7_3_W0_data = W0_data[31:24];
  assign mem_7_3_W0_en = W0_en & W0_addr_sel == 8'h7;
  assign mem_7_3_W0_mask = W0_mask[3];
  assign mem_7_4_R0_addr = R0_addr[25:0];
  assign mem_7_4_R0_clk = R0_clk;
  assign mem_7_4_R0_en = R0_en & R0_addr_sel == 8'h7;
  assign mem_7_4_W0_addr = W0_addr[25:0];
  assign mem_7_4_W0_clk = W0_clk;
  assign mem_7_4_W0_data = W0_data[39:32];
  assign mem_7_4_W0_en = W0_en & W0_addr_sel == 8'h7;
  assign mem_7_4_W0_mask = W0_mask[4];
  assign mem_7_5_R0_addr = R0_addr[25:0];
  assign mem_7_5_R0_clk = R0_clk;
  assign mem_7_5_R0_en = R0_en & R0_addr_sel == 8'h7;
  assign mem_7_5_W0_addr = W0_addr[25:0];
  assign mem_7_5_W0_clk = W0_clk;
  assign mem_7_5_W0_data = W0_data[47:40];
  assign mem_7_5_W0_en = W0_en & W0_addr_sel == 8'h7;
  assign mem_7_5_W0_mask = W0_mask[5];
  assign mem_7_6_R0_addr = R0_addr[25:0];
  assign mem_7_6_R0_clk = R0_clk;
  assign mem_7_6_R0_en = R0_en & R0_addr_sel == 8'h7;
  assign mem_7_6_W0_addr = W0_addr[25:0];
  assign mem_7_6_W0_clk = W0_clk;
  assign mem_7_6_W0_data = W0_data[55:48];
  assign mem_7_6_W0_en = W0_en & W0_addr_sel == 8'h7;
  assign mem_7_6_W0_mask = W0_mask[6];
  assign mem_7_7_R0_addr = R0_addr[25:0];
  assign mem_7_7_R0_clk = R0_clk;
  assign mem_7_7_R0_en = R0_en & R0_addr_sel == 8'h7;
  assign mem_7_7_W0_addr = W0_addr[25:0];
  assign mem_7_7_W0_clk = W0_clk;
  assign mem_7_7_W0_data = W0_data[63:56];
  assign mem_7_7_W0_en = W0_en & W0_addr_sel == 8'h7;
  assign mem_7_7_W0_mask = W0_mask[7];
  assign mem_8_0_R0_addr = R0_addr[25:0];
  assign mem_8_0_R0_clk = R0_clk;
  assign mem_8_0_R0_en = R0_en & R0_addr_sel == 8'h8;
  assign mem_8_0_W0_addr = W0_addr[25:0];
  assign mem_8_0_W0_clk = W0_clk;
  assign mem_8_0_W0_data = W0_data[7:0];
  assign mem_8_0_W0_en = W0_en & W0_addr_sel == 8'h8;
  assign mem_8_0_W0_mask = W0_mask[0];
  assign mem_8_1_R0_addr = R0_addr[25:0];
  assign mem_8_1_R0_clk = R0_clk;
  assign mem_8_1_R0_en = R0_en & R0_addr_sel == 8'h8;
  assign mem_8_1_W0_addr = W0_addr[25:0];
  assign mem_8_1_W0_clk = W0_clk;
  assign mem_8_1_W0_data = W0_data[15:8];
  assign mem_8_1_W0_en = W0_en & W0_addr_sel == 8'h8;
  assign mem_8_1_W0_mask = W0_mask[1];
  assign mem_8_2_R0_addr = R0_addr[25:0];
  assign mem_8_2_R0_clk = R0_clk;
  assign mem_8_2_R0_en = R0_en & R0_addr_sel == 8'h8;
  assign mem_8_2_W0_addr = W0_addr[25:0];
  assign mem_8_2_W0_clk = W0_clk;
  assign mem_8_2_W0_data = W0_data[23:16];
  assign mem_8_2_W0_en = W0_en & W0_addr_sel == 8'h8;
  assign mem_8_2_W0_mask = W0_mask[2];
  assign mem_8_3_R0_addr = R0_addr[25:0];
  assign mem_8_3_R0_clk = R0_clk;
  assign mem_8_3_R0_en = R0_en & R0_addr_sel == 8'h8;
  assign mem_8_3_W0_addr = W0_addr[25:0];
  assign mem_8_3_W0_clk = W0_clk;
  assign mem_8_3_W0_data = W0_data[31:24];
  assign mem_8_3_W0_en = W0_en & W0_addr_sel == 8'h8;
  assign mem_8_3_W0_mask = W0_mask[3];
  assign mem_8_4_R0_addr = R0_addr[25:0];
  assign mem_8_4_R0_clk = R0_clk;
  assign mem_8_4_R0_en = R0_en & R0_addr_sel == 8'h8;
  assign mem_8_4_W0_addr = W0_addr[25:0];
  assign mem_8_4_W0_clk = W0_clk;
  assign mem_8_4_W0_data = W0_data[39:32];
  assign mem_8_4_W0_en = W0_en & W0_addr_sel == 8'h8;
  assign mem_8_4_W0_mask = W0_mask[4];
  assign mem_8_5_R0_addr = R0_addr[25:0];
  assign mem_8_5_R0_clk = R0_clk;
  assign mem_8_5_R0_en = R0_en & R0_addr_sel == 8'h8;
  assign mem_8_5_W0_addr = W0_addr[25:0];
  assign mem_8_5_W0_clk = W0_clk;
  assign mem_8_5_W0_data = W0_data[47:40];
  assign mem_8_5_W0_en = W0_en & W0_addr_sel == 8'h8;
  assign mem_8_5_W0_mask = W0_mask[5];
  assign mem_8_6_R0_addr = R0_addr[25:0];
  assign mem_8_6_R0_clk = R0_clk;
  assign mem_8_6_R0_en = R0_en & R0_addr_sel == 8'h8;
  assign mem_8_6_W0_addr = W0_addr[25:0];
  assign mem_8_6_W0_clk = W0_clk;
  assign mem_8_6_W0_data = W0_data[55:48];
  assign mem_8_6_W0_en = W0_en & W0_addr_sel == 8'h8;
  assign mem_8_6_W0_mask = W0_mask[6];
  assign mem_8_7_R0_addr = R0_addr[25:0];
  assign mem_8_7_R0_clk = R0_clk;
  assign mem_8_7_R0_en = R0_en & R0_addr_sel == 8'h8;
  assign mem_8_7_W0_addr = W0_addr[25:0];
  assign mem_8_7_W0_clk = W0_clk;
  assign mem_8_7_W0_data = W0_data[63:56];
  assign mem_8_7_W0_en = W0_en & W0_addr_sel == 8'h8;
  assign mem_8_7_W0_mask = W0_mask[7];
  assign mem_9_0_R0_addr = R0_addr[25:0];
  assign mem_9_0_R0_clk = R0_clk;
  assign mem_9_0_R0_en = R0_en & R0_addr_sel == 8'h9;
  assign mem_9_0_W0_addr = W0_addr[25:0];
  assign mem_9_0_W0_clk = W0_clk;
  assign mem_9_0_W0_data = W0_data[7:0];
  assign mem_9_0_W0_en = W0_en & W0_addr_sel == 8'h9;
  assign mem_9_0_W0_mask = W0_mask[0];
  assign mem_9_1_R0_addr = R0_addr[25:0];
  assign mem_9_1_R0_clk = R0_clk;
  assign mem_9_1_R0_en = R0_en & R0_addr_sel == 8'h9;
  assign mem_9_1_W0_addr = W0_addr[25:0];
  assign mem_9_1_W0_clk = W0_clk;
  assign mem_9_1_W0_data = W0_data[15:8];
  assign mem_9_1_W0_en = W0_en & W0_addr_sel == 8'h9;
  assign mem_9_1_W0_mask = W0_mask[1];
  assign mem_9_2_R0_addr = R0_addr[25:0];
  assign mem_9_2_R0_clk = R0_clk;
  assign mem_9_2_R0_en = R0_en & R0_addr_sel == 8'h9;
  assign mem_9_2_W0_addr = W0_addr[25:0];
  assign mem_9_2_W0_clk = W0_clk;
  assign mem_9_2_W0_data = W0_data[23:16];
  assign mem_9_2_W0_en = W0_en & W0_addr_sel == 8'h9;
  assign mem_9_2_W0_mask = W0_mask[2];
  assign mem_9_3_R0_addr = R0_addr[25:0];
  assign mem_9_3_R0_clk = R0_clk;
  assign mem_9_3_R0_en = R0_en & R0_addr_sel == 8'h9;
  assign mem_9_3_W0_addr = W0_addr[25:0];
  assign mem_9_3_W0_clk = W0_clk;
  assign mem_9_3_W0_data = W0_data[31:24];
  assign mem_9_3_W0_en = W0_en & W0_addr_sel == 8'h9;
  assign mem_9_3_W0_mask = W0_mask[3];
  assign mem_9_4_R0_addr = R0_addr[25:0];
  assign mem_9_4_R0_clk = R0_clk;
  assign mem_9_4_R0_en = R0_en & R0_addr_sel == 8'h9;
  assign mem_9_4_W0_addr = W0_addr[25:0];
  assign mem_9_4_W0_clk = W0_clk;
  assign mem_9_4_W0_data = W0_data[39:32];
  assign mem_9_4_W0_en = W0_en & W0_addr_sel == 8'h9;
  assign mem_9_4_W0_mask = W0_mask[4];
  assign mem_9_5_R0_addr = R0_addr[25:0];
  assign mem_9_5_R0_clk = R0_clk;
  assign mem_9_5_R0_en = R0_en & R0_addr_sel == 8'h9;
  assign mem_9_5_W0_addr = W0_addr[25:0];
  assign mem_9_5_W0_clk = W0_clk;
  assign mem_9_5_W0_data = W0_data[47:40];
  assign mem_9_5_W0_en = W0_en & W0_addr_sel == 8'h9;
  assign mem_9_5_W0_mask = W0_mask[5];
  assign mem_9_6_R0_addr = R0_addr[25:0];
  assign mem_9_6_R0_clk = R0_clk;
  assign mem_9_6_R0_en = R0_en & R0_addr_sel == 8'h9;
  assign mem_9_6_W0_addr = W0_addr[25:0];
  assign mem_9_6_W0_clk = W0_clk;
  assign mem_9_6_W0_data = W0_data[55:48];
  assign mem_9_6_W0_en = W0_en & W0_addr_sel == 8'h9;
  assign mem_9_6_W0_mask = W0_mask[6];
  assign mem_9_7_R0_addr = R0_addr[25:0];
  assign mem_9_7_R0_clk = R0_clk;
  assign mem_9_7_R0_en = R0_en & R0_addr_sel == 8'h9;
  assign mem_9_7_W0_addr = W0_addr[25:0];
  assign mem_9_7_W0_clk = W0_clk;
  assign mem_9_7_W0_data = W0_data[63:56];
  assign mem_9_7_W0_en = W0_en & W0_addr_sel == 8'h9;
  assign mem_9_7_W0_mask = W0_mask[7];
  assign mem_10_0_R0_addr = R0_addr[25:0];
  assign mem_10_0_R0_clk = R0_clk;
  assign mem_10_0_R0_en = R0_en & R0_addr_sel == 8'ha;
  assign mem_10_0_W0_addr = W0_addr[25:0];
  assign mem_10_0_W0_clk = W0_clk;
  assign mem_10_0_W0_data = W0_data[7:0];
  assign mem_10_0_W0_en = W0_en & W0_addr_sel == 8'ha;
  assign mem_10_0_W0_mask = W0_mask[0];
  assign mem_10_1_R0_addr = R0_addr[25:0];
  assign mem_10_1_R0_clk = R0_clk;
  assign mem_10_1_R0_en = R0_en & R0_addr_sel == 8'ha;
  assign mem_10_1_W0_addr = W0_addr[25:0];
  assign mem_10_1_W0_clk = W0_clk;
  assign mem_10_1_W0_data = W0_data[15:8];
  assign mem_10_1_W0_en = W0_en & W0_addr_sel == 8'ha;
  assign mem_10_1_W0_mask = W0_mask[1];
  assign mem_10_2_R0_addr = R0_addr[25:0];
  assign mem_10_2_R0_clk = R0_clk;
  assign mem_10_2_R0_en = R0_en & R0_addr_sel == 8'ha;
  assign mem_10_2_W0_addr = W0_addr[25:0];
  assign mem_10_2_W0_clk = W0_clk;
  assign mem_10_2_W0_data = W0_data[23:16];
  assign mem_10_2_W0_en = W0_en & W0_addr_sel == 8'ha;
  assign mem_10_2_W0_mask = W0_mask[2];
  assign mem_10_3_R0_addr = R0_addr[25:0];
  assign mem_10_3_R0_clk = R0_clk;
  assign mem_10_3_R0_en = R0_en & R0_addr_sel == 8'ha;
  assign mem_10_3_W0_addr = W0_addr[25:0];
  assign mem_10_3_W0_clk = W0_clk;
  assign mem_10_3_W0_data = W0_data[31:24];
  assign mem_10_3_W0_en = W0_en & W0_addr_sel == 8'ha;
  assign mem_10_3_W0_mask = W0_mask[3];
  assign mem_10_4_R0_addr = R0_addr[25:0];
  assign mem_10_4_R0_clk = R0_clk;
  assign mem_10_4_R0_en = R0_en & R0_addr_sel == 8'ha;
  assign mem_10_4_W0_addr = W0_addr[25:0];
  assign mem_10_4_W0_clk = W0_clk;
  assign mem_10_4_W0_data = W0_data[39:32];
  assign mem_10_4_W0_en = W0_en & W0_addr_sel == 8'ha;
  assign mem_10_4_W0_mask = W0_mask[4];
  assign mem_10_5_R0_addr = R0_addr[25:0];
  assign mem_10_5_R0_clk = R0_clk;
  assign mem_10_5_R0_en = R0_en & R0_addr_sel == 8'ha;
  assign mem_10_5_W0_addr = W0_addr[25:0];
  assign mem_10_5_W0_clk = W0_clk;
  assign mem_10_5_W0_data = W0_data[47:40];
  assign mem_10_5_W0_en = W0_en & W0_addr_sel == 8'ha;
  assign mem_10_5_W0_mask = W0_mask[5];
  assign mem_10_6_R0_addr = R0_addr[25:0];
  assign mem_10_6_R0_clk = R0_clk;
  assign mem_10_6_R0_en = R0_en & R0_addr_sel == 8'ha;
  assign mem_10_6_W0_addr = W0_addr[25:0];
  assign mem_10_6_W0_clk = W0_clk;
  assign mem_10_6_W0_data = W0_data[55:48];
  assign mem_10_6_W0_en = W0_en & W0_addr_sel == 8'ha;
  assign mem_10_6_W0_mask = W0_mask[6];
  assign mem_10_7_R0_addr = R0_addr[25:0];
  assign mem_10_7_R0_clk = R0_clk;
  assign mem_10_7_R0_en = R0_en & R0_addr_sel == 8'ha;
  assign mem_10_7_W0_addr = W0_addr[25:0];
  assign mem_10_7_W0_clk = W0_clk;
  assign mem_10_7_W0_data = W0_data[63:56];
  assign mem_10_7_W0_en = W0_en & W0_addr_sel == 8'ha;
  assign mem_10_7_W0_mask = W0_mask[7];
  assign mem_11_0_R0_addr = R0_addr[25:0];
  assign mem_11_0_R0_clk = R0_clk;
  assign mem_11_0_R0_en = R0_en & R0_addr_sel == 8'hb;
  assign mem_11_0_W0_addr = W0_addr[25:0];
  assign mem_11_0_W0_clk = W0_clk;
  assign mem_11_0_W0_data = W0_data[7:0];
  assign mem_11_0_W0_en = W0_en & W0_addr_sel == 8'hb;
  assign mem_11_0_W0_mask = W0_mask[0];
  assign mem_11_1_R0_addr = R0_addr[25:0];
  assign mem_11_1_R0_clk = R0_clk;
  assign mem_11_1_R0_en = R0_en & R0_addr_sel == 8'hb;
  assign mem_11_1_W0_addr = W0_addr[25:0];
  assign mem_11_1_W0_clk = W0_clk;
  assign mem_11_1_W0_data = W0_data[15:8];
  assign mem_11_1_W0_en = W0_en & W0_addr_sel == 8'hb;
  assign mem_11_1_W0_mask = W0_mask[1];
  assign mem_11_2_R0_addr = R0_addr[25:0];
  assign mem_11_2_R0_clk = R0_clk;
  assign mem_11_2_R0_en = R0_en & R0_addr_sel == 8'hb;
  assign mem_11_2_W0_addr = W0_addr[25:0];
  assign mem_11_2_W0_clk = W0_clk;
  assign mem_11_2_W0_data = W0_data[23:16];
  assign mem_11_2_W0_en = W0_en & W0_addr_sel == 8'hb;
  assign mem_11_2_W0_mask = W0_mask[2];
  assign mem_11_3_R0_addr = R0_addr[25:0];
  assign mem_11_3_R0_clk = R0_clk;
  assign mem_11_3_R0_en = R0_en & R0_addr_sel == 8'hb;
  assign mem_11_3_W0_addr = W0_addr[25:0];
  assign mem_11_3_W0_clk = W0_clk;
  assign mem_11_3_W0_data = W0_data[31:24];
  assign mem_11_3_W0_en = W0_en & W0_addr_sel == 8'hb;
  assign mem_11_3_W0_mask = W0_mask[3];
  assign mem_11_4_R0_addr = R0_addr[25:0];
  assign mem_11_4_R0_clk = R0_clk;
  assign mem_11_4_R0_en = R0_en & R0_addr_sel == 8'hb;
  assign mem_11_4_W0_addr = W0_addr[25:0];
  assign mem_11_4_W0_clk = W0_clk;
  assign mem_11_4_W0_data = W0_data[39:32];
  assign mem_11_4_W0_en = W0_en & W0_addr_sel == 8'hb;
  assign mem_11_4_W0_mask = W0_mask[4];
  assign mem_11_5_R0_addr = R0_addr[25:0];
  assign mem_11_5_R0_clk = R0_clk;
  assign mem_11_5_R0_en = R0_en & R0_addr_sel == 8'hb;
  assign mem_11_5_W0_addr = W0_addr[25:0];
  assign mem_11_5_W0_clk = W0_clk;
  assign mem_11_5_W0_data = W0_data[47:40];
  assign mem_11_5_W0_en = W0_en & W0_addr_sel == 8'hb;
  assign mem_11_5_W0_mask = W0_mask[5];
  assign mem_11_6_R0_addr = R0_addr[25:0];
  assign mem_11_6_R0_clk = R0_clk;
  assign mem_11_6_R0_en = R0_en & R0_addr_sel == 8'hb;
  assign mem_11_6_W0_addr = W0_addr[25:0];
  assign mem_11_6_W0_clk = W0_clk;
  assign mem_11_6_W0_data = W0_data[55:48];
  assign mem_11_6_W0_en = W0_en & W0_addr_sel == 8'hb;
  assign mem_11_6_W0_mask = W0_mask[6];
  assign mem_11_7_R0_addr = R0_addr[25:0];
  assign mem_11_7_R0_clk = R0_clk;
  assign mem_11_7_R0_en = R0_en & R0_addr_sel == 8'hb;
  assign mem_11_7_W0_addr = W0_addr[25:0];
  assign mem_11_7_W0_clk = W0_clk;
  assign mem_11_7_W0_data = W0_data[63:56];
  assign mem_11_7_W0_en = W0_en & W0_addr_sel == 8'hb;
  assign mem_11_7_W0_mask = W0_mask[7];
  assign mem_12_0_R0_addr = R0_addr[25:0];
  assign mem_12_0_R0_clk = R0_clk;
  assign mem_12_0_R0_en = R0_en & R0_addr_sel == 8'hc;
  assign mem_12_0_W0_addr = W0_addr[25:0];
  assign mem_12_0_W0_clk = W0_clk;
  assign mem_12_0_W0_data = W0_data[7:0];
  assign mem_12_0_W0_en = W0_en & W0_addr_sel == 8'hc;
  assign mem_12_0_W0_mask = W0_mask[0];
  assign mem_12_1_R0_addr = R0_addr[25:0];
  assign mem_12_1_R0_clk = R0_clk;
  assign mem_12_1_R0_en = R0_en & R0_addr_sel == 8'hc;
  assign mem_12_1_W0_addr = W0_addr[25:0];
  assign mem_12_1_W0_clk = W0_clk;
  assign mem_12_1_W0_data = W0_data[15:8];
  assign mem_12_1_W0_en = W0_en & W0_addr_sel == 8'hc;
  assign mem_12_1_W0_mask = W0_mask[1];
  assign mem_12_2_R0_addr = R0_addr[25:0];
  assign mem_12_2_R0_clk = R0_clk;
  assign mem_12_2_R0_en = R0_en & R0_addr_sel == 8'hc;
  assign mem_12_2_W0_addr = W0_addr[25:0];
  assign mem_12_2_W0_clk = W0_clk;
  assign mem_12_2_W0_data = W0_data[23:16];
  assign mem_12_2_W0_en = W0_en & W0_addr_sel == 8'hc;
  assign mem_12_2_W0_mask = W0_mask[2];
  assign mem_12_3_R0_addr = R0_addr[25:0];
  assign mem_12_3_R0_clk = R0_clk;
  assign mem_12_3_R0_en = R0_en & R0_addr_sel == 8'hc;
  assign mem_12_3_W0_addr = W0_addr[25:0];
  assign mem_12_3_W0_clk = W0_clk;
  assign mem_12_3_W0_data = W0_data[31:24];
  assign mem_12_3_W0_en = W0_en & W0_addr_sel == 8'hc;
  assign mem_12_3_W0_mask = W0_mask[3];
  assign mem_12_4_R0_addr = R0_addr[25:0];
  assign mem_12_4_R0_clk = R0_clk;
  assign mem_12_4_R0_en = R0_en & R0_addr_sel == 8'hc;
  assign mem_12_4_W0_addr = W0_addr[25:0];
  assign mem_12_4_W0_clk = W0_clk;
  assign mem_12_4_W0_data = W0_data[39:32];
  assign mem_12_4_W0_en = W0_en & W0_addr_sel == 8'hc;
  assign mem_12_4_W0_mask = W0_mask[4];
  assign mem_12_5_R0_addr = R0_addr[25:0];
  assign mem_12_5_R0_clk = R0_clk;
  assign mem_12_5_R0_en = R0_en & R0_addr_sel == 8'hc;
  assign mem_12_5_W0_addr = W0_addr[25:0];
  assign mem_12_5_W0_clk = W0_clk;
  assign mem_12_5_W0_data = W0_data[47:40];
  assign mem_12_5_W0_en = W0_en & W0_addr_sel == 8'hc;
  assign mem_12_5_W0_mask = W0_mask[5];
  assign mem_12_6_R0_addr = R0_addr[25:0];
  assign mem_12_6_R0_clk = R0_clk;
  assign mem_12_6_R0_en = R0_en & R0_addr_sel == 8'hc;
  assign mem_12_6_W0_addr = W0_addr[25:0];
  assign mem_12_6_W0_clk = W0_clk;
  assign mem_12_6_W0_data = W0_data[55:48];
  assign mem_12_6_W0_en = W0_en & W0_addr_sel == 8'hc;
  assign mem_12_6_W0_mask = W0_mask[6];
  assign mem_12_7_R0_addr = R0_addr[25:0];
  assign mem_12_7_R0_clk = R0_clk;
  assign mem_12_7_R0_en = R0_en & R0_addr_sel == 8'hc;
  assign mem_12_7_W0_addr = W0_addr[25:0];
  assign mem_12_7_W0_clk = W0_clk;
  assign mem_12_7_W0_data = W0_data[63:56];
  assign mem_12_7_W0_en = W0_en & W0_addr_sel == 8'hc;
  assign mem_12_7_W0_mask = W0_mask[7];
  assign mem_13_0_R0_addr = R0_addr[25:0];
  assign mem_13_0_R0_clk = R0_clk;
  assign mem_13_0_R0_en = R0_en & R0_addr_sel == 8'hd;
  assign mem_13_0_W0_addr = W0_addr[25:0];
  assign mem_13_0_W0_clk = W0_clk;
  assign mem_13_0_W0_data = W0_data[7:0];
  assign mem_13_0_W0_en = W0_en & W0_addr_sel == 8'hd;
  assign mem_13_0_W0_mask = W0_mask[0];
  assign mem_13_1_R0_addr = R0_addr[25:0];
  assign mem_13_1_R0_clk = R0_clk;
  assign mem_13_1_R0_en = R0_en & R0_addr_sel == 8'hd;
  assign mem_13_1_W0_addr = W0_addr[25:0];
  assign mem_13_1_W0_clk = W0_clk;
  assign mem_13_1_W0_data = W0_data[15:8];
  assign mem_13_1_W0_en = W0_en & W0_addr_sel == 8'hd;
  assign mem_13_1_W0_mask = W0_mask[1];
  assign mem_13_2_R0_addr = R0_addr[25:0];
  assign mem_13_2_R0_clk = R0_clk;
  assign mem_13_2_R0_en = R0_en & R0_addr_sel == 8'hd;
  assign mem_13_2_W0_addr = W0_addr[25:0];
  assign mem_13_2_W0_clk = W0_clk;
  assign mem_13_2_W0_data = W0_data[23:16];
  assign mem_13_2_W0_en = W0_en & W0_addr_sel == 8'hd;
  assign mem_13_2_W0_mask = W0_mask[2];
  assign mem_13_3_R0_addr = R0_addr[25:0];
  assign mem_13_3_R0_clk = R0_clk;
  assign mem_13_3_R0_en = R0_en & R0_addr_sel == 8'hd;
  assign mem_13_3_W0_addr = W0_addr[25:0];
  assign mem_13_3_W0_clk = W0_clk;
  assign mem_13_3_W0_data = W0_data[31:24];
  assign mem_13_3_W0_en = W0_en & W0_addr_sel == 8'hd;
  assign mem_13_3_W0_mask = W0_mask[3];
  assign mem_13_4_R0_addr = R0_addr[25:0];
  assign mem_13_4_R0_clk = R0_clk;
  assign mem_13_4_R0_en = R0_en & R0_addr_sel == 8'hd;
  assign mem_13_4_W0_addr = W0_addr[25:0];
  assign mem_13_4_W0_clk = W0_clk;
  assign mem_13_4_W0_data = W0_data[39:32];
  assign mem_13_4_W0_en = W0_en & W0_addr_sel == 8'hd;
  assign mem_13_4_W0_mask = W0_mask[4];
  assign mem_13_5_R0_addr = R0_addr[25:0];
  assign mem_13_5_R0_clk = R0_clk;
  assign mem_13_5_R0_en = R0_en & R0_addr_sel == 8'hd;
  assign mem_13_5_W0_addr = W0_addr[25:0];
  assign mem_13_5_W0_clk = W0_clk;
  assign mem_13_5_W0_data = W0_data[47:40];
  assign mem_13_5_W0_en = W0_en & W0_addr_sel == 8'hd;
  assign mem_13_5_W0_mask = W0_mask[5];
  assign mem_13_6_R0_addr = R0_addr[25:0];
  assign mem_13_6_R0_clk = R0_clk;
  assign mem_13_6_R0_en = R0_en & R0_addr_sel == 8'hd;
  assign mem_13_6_W0_addr = W0_addr[25:0];
  assign mem_13_6_W0_clk = W0_clk;
  assign mem_13_6_W0_data = W0_data[55:48];
  assign mem_13_6_W0_en = W0_en & W0_addr_sel == 8'hd;
  assign mem_13_6_W0_mask = W0_mask[6];
  assign mem_13_7_R0_addr = R0_addr[25:0];
  assign mem_13_7_R0_clk = R0_clk;
  assign mem_13_7_R0_en = R0_en & R0_addr_sel == 8'hd;
  assign mem_13_7_W0_addr = W0_addr[25:0];
  assign mem_13_7_W0_clk = W0_clk;
  assign mem_13_7_W0_data = W0_data[63:56];
  assign mem_13_7_W0_en = W0_en & W0_addr_sel == 8'hd;
  assign mem_13_7_W0_mask = W0_mask[7];
  assign mem_14_0_R0_addr = R0_addr[25:0];
  assign mem_14_0_R0_clk = R0_clk;
  assign mem_14_0_R0_en = R0_en & R0_addr_sel == 8'he;
  assign mem_14_0_W0_addr = W0_addr[25:0];
  assign mem_14_0_W0_clk = W0_clk;
  assign mem_14_0_W0_data = W0_data[7:0];
  assign mem_14_0_W0_en = W0_en & W0_addr_sel == 8'he;
  assign mem_14_0_W0_mask = W0_mask[0];
  assign mem_14_1_R0_addr = R0_addr[25:0];
  assign mem_14_1_R0_clk = R0_clk;
  assign mem_14_1_R0_en = R0_en & R0_addr_sel == 8'he;
  assign mem_14_1_W0_addr = W0_addr[25:0];
  assign mem_14_1_W0_clk = W0_clk;
  assign mem_14_1_W0_data = W0_data[15:8];
  assign mem_14_1_W0_en = W0_en & W0_addr_sel == 8'he;
  assign mem_14_1_W0_mask = W0_mask[1];
  assign mem_14_2_R0_addr = R0_addr[25:0];
  assign mem_14_2_R0_clk = R0_clk;
  assign mem_14_2_R0_en = R0_en & R0_addr_sel == 8'he;
  assign mem_14_2_W0_addr = W0_addr[25:0];
  assign mem_14_2_W0_clk = W0_clk;
  assign mem_14_2_W0_data = W0_data[23:16];
  assign mem_14_2_W0_en = W0_en & W0_addr_sel == 8'he;
  assign mem_14_2_W0_mask = W0_mask[2];
  assign mem_14_3_R0_addr = R0_addr[25:0];
  assign mem_14_3_R0_clk = R0_clk;
  assign mem_14_3_R0_en = R0_en & R0_addr_sel == 8'he;
  assign mem_14_3_W0_addr = W0_addr[25:0];
  assign mem_14_3_W0_clk = W0_clk;
  assign mem_14_3_W0_data = W0_data[31:24];
  assign mem_14_3_W0_en = W0_en & W0_addr_sel == 8'he;
  assign mem_14_3_W0_mask = W0_mask[3];
  assign mem_14_4_R0_addr = R0_addr[25:0];
  assign mem_14_4_R0_clk = R0_clk;
  assign mem_14_4_R0_en = R0_en & R0_addr_sel == 8'he;
  assign mem_14_4_W0_addr = W0_addr[25:0];
  assign mem_14_4_W0_clk = W0_clk;
  assign mem_14_4_W0_data = W0_data[39:32];
  assign mem_14_4_W0_en = W0_en & W0_addr_sel == 8'he;
  assign mem_14_4_W0_mask = W0_mask[4];
  assign mem_14_5_R0_addr = R0_addr[25:0];
  assign mem_14_5_R0_clk = R0_clk;
  assign mem_14_5_R0_en = R0_en & R0_addr_sel == 8'he;
  assign mem_14_5_W0_addr = W0_addr[25:0];
  assign mem_14_5_W0_clk = W0_clk;
  assign mem_14_5_W0_data = W0_data[47:40];
  assign mem_14_5_W0_en = W0_en & W0_addr_sel == 8'he;
  assign mem_14_5_W0_mask = W0_mask[5];
  assign mem_14_6_R0_addr = R0_addr[25:0];
  assign mem_14_6_R0_clk = R0_clk;
  assign mem_14_6_R0_en = R0_en & R0_addr_sel == 8'he;
  assign mem_14_6_W0_addr = W0_addr[25:0];
  assign mem_14_6_W0_clk = W0_clk;
  assign mem_14_6_W0_data = W0_data[55:48];
  assign mem_14_6_W0_en = W0_en & W0_addr_sel == 8'he;
  assign mem_14_6_W0_mask = W0_mask[6];
  assign mem_14_7_R0_addr = R0_addr[25:0];
  assign mem_14_7_R0_clk = R0_clk;
  assign mem_14_7_R0_en = R0_en & R0_addr_sel == 8'he;
  assign mem_14_7_W0_addr = W0_addr[25:0];
  assign mem_14_7_W0_clk = W0_clk;
  assign mem_14_7_W0_data = W0_data[63:56];
  assign mem_14_7_W0_en = W0_en & W0_addr_sel == 8'he;
  assign mem_14_7_W0_mask = W0_mask[7];
  assign mem_15_0_R0_addr = R0_addr[25:0];
  assign mem_15_0_R0_clk = R0_clk;
  assign mem_15_0_R0_en = R0_en & R0_addr_sel == 8'hf;
  assign mem_15_0_W0_addr = W0_addr[25:0];
  assign mem_15_0_W0_clk = W0_clk;
  assign mem_15_0_W0_data = W0_data[7:0];
  assign mem_15_0_W0_en = W0_en & W0_addr_sel == 8'hf;
  assign mem_15_0_W0_mask = W0_mask[0];
  assign mem_15_1_R0_addr = R0_addr[25:0];
  assign mem_15_1_R0_clk = R0_clk;
  assign mem_15_1_R0_en = R0_en & R0_addr_sel == 8'hf;
  assign mem_15_1_W0_addr = W0_addr[25:0];
  assign mem_15_1_W0_clk = W0_clk;
  assign mem_15_1_W0_data = W0_data[15:8];
  assign mem_15_1_W0_en = W0_en & W0_addr_sel == 8'hf;
  assign mem_15_1_W0_mask = W0_mask[1];
  assign mem_15_2_R0_addr = R0_addr[25:0];
  assign mem_15_2_R0_clk = R0_clk;
  assign mem_15_2_R0_en = R0_en & R0_addr_sel == 8'hf;
  assign mem_15_2_W0_addr = W0_addr[25:0];
  assign mem_15_2_W0_clk = W0_clk;
  assign mem_15_2_W0_data = W0_data[23:16];
  assign mem_15_2_W0_en = W0_en & W0_addr_sel == 8'hf;
  assign mem_15_2_W0_mask = W0_mask[2];
  assign mem_15_3_R0_addr = R0_addr[25:0];
  assign mem_15_3_R0_clk = R0_clk;
  assign mem_15_3_R0_en = R0_en & R0_addr_sel == 8'hf;
  assign mem_15_3_W0_addr = W0_addr[25:0];
  assign mem_15_3_W0_clk = W0_clk;
  assign mem_15_3_W0_data = W0_data[31:24];
  assign mem_15_3_W0_en = W0_en & W0_addr_sel == 8'hf;
  assign mem_15_3_W0_mask = W0_mask[3];
  assign mem_15_4_R0_addr = R0_addr[25:0];
  assign mem_15_4_R0_clk = R0_clk;
  assign mem_15_4_R0_en = R0_en & R0_addr_sel == 8'hf;
  assign mem_15_4_W0_addr = W0_addr[25:0];
  assign mem_15_4_W0_clk = W0_clk;
  assign mem_15_4_W0_data = W0_data[39:32];
  assign mem_15_4_W0_en = W0_en & W0_addr_sel == 8'hf;
  assign mem_15_4_W0_mask = W0_mask[4];
  assign mem_15_5_R0_addr = R0_addr[25:0];
  assign mem_15_5_R0_clk = R0_clk;
  assign mem_15_5_R0_en = R0_en & R0_addr_sel == 8'hf;
  assign mem_15_5_W0_addr = W0_addr[25:0];
  assign mem_15_5_W0_clk = W0_clk;
  assign mem_15_5_W0_data = W0_data[47:40];
  assign mem_15_5_W0_en = W0_en & W0_addr_sel == 8'hf;
  assign mem_15_5_W0_mask = W0_mask[5];
  assign mem_15_6_R0_addr = R0_addr[25:0];
  assign mem_15_6_R0_clk = R0_clk;
  assign mem_15_6_R0_en = R0_en & R0_addr_sel == 8'hf;
  assign mem_15_6_W0_addr = W0_addr[25:0];
  assign mem_15_6_W0_clk = W0_clk;
  assign mem_15_6_W0_data = W0_data[55:48];
  assign mem_15_6_W0_en = W0_en & W0_addr_sel == 8'hf;
  assign mem_15_6_W0_mask = W0_mask[6];
  assign mem_15_7_R0_addr = R0_addr[25:0];
  assign mem_15_7_R0_clk = R0_clk;
  assign mem_15_7_R0_en = R0_en & R0_addr_sel == 8'hf;
  assign mem_15_7_W0_addr = W0_addr[25:0];
  assign mem_15_7_W0_clk = W0_clk;
  assign mem_15_7_W0_data = W0_data[63:56];
  assign mem_15_7_W0_en = W0_en & W0_addr_sel == 8'hf;
  assign mem_15_7_W0_mask = W0_mask[7];
  assign mem_16_0_R0_addr = R0_addr[25:0];
  assign mem_16_0_R0_clk = R0_clk;
  assign mem_16_0_R0_en = R0_en & R0_addr_sel == 8'h10;
  assign mem_16_0_W0_addr = W0_addr[25:0];
  assign mem_16_0_W0_clk = W0_clk;
  assign mem_16_0_W0_data = W0_data[7:0];
  assign mem_16_0_W0_en = W0_en & W0_addr_sel == 8'h10;
  assign mem_16_0_W0_mask = W0_mask[0];
  assign mem_16_1_R0_addr = R0_addr[25:0];
  assign mem_16_1_R0_clk = R0_clk;
  assign mem_16_1_R0_en = R0_en & R0_addr_sel == 8'h10;
  assign mem_16_1_W0_addr = W0_addr[25:0];
  assign mem_16_1_W0_clk = W0_clk;
  assign mem_16_1_W0_data = W0_data[15:8];
  assign mem_16_1_W0_en = W0_en & W0_addr_sel == 8'h10;
  assign mem_16_1_W0_mask = W0_mask[1];
  assign mem_16_2_R0_addr = R0_addr[25:0];
  assign mem_16_2_R0_clk = R0_clk;
  assign mem_16_2_R0_en = R0_en & R0_addr_sel == 8'h10;
  assign mem_16_2_W0_addr = W0_addr[25:0];
  assign mem_16_2_W0_clk = W0_clk;
  assign mem_16_2_W0_data = W0_data[23:16];
  assign mem_16_2_W0_en = W0_en & W0_addr_sel == 8'h10;
  assign mem_16_2_W0_mask = W0_mask[2];
  assign mem_16_3_R0_addr = R0_addr[25:0];
  assign mem_16_3_R0_clk = R0_clk;
  assign mem_16_3_R0_en = R0_en & R0_addr_sel == 8'h10;
  assign mem_16_3_W0_addr = W0_addr[25:0];
  assign mem_16_3_W0_clk = W0_clk;
  assign mem_16_3_W0_data = W0_data[31:24];
  assign mem_16_3_W0_en = W0_en & W0_addr_sel == 8'h10;
  assign mem_16_3_W0_mask = W0_mask[3];
  assign mem_16_4_R0_addr = R0_addr[25:0];
  assign mem_16_4_R0_clk = R0_clk;
  assign mem_16_4_R0_en = R0_en & R0_addr_sel == 8'h10;
  assign mem_16_4_W0_addr = W0_addr[25:0];
  assign mem_16_4_W0_clk = W0_clk;
  assign mem_16_4_W0_data = W0_data[39:32];
  assign mem_16_4_W0_en = W0_en & W0_addr_sel == 8'h10;
  assign mem_16_4_W0_mask = W0_mask[4];
  assign mem_16_5_R0_addr = R0_addr[25:0];
  assign mem_16_5_R0_clk = R0_clk;
  assign mem_16_5_R0_en = R0_en & R0_addr_sel == 8'h10;
  assign mem_16_5_W0_addr = W0_addr[25:0];
  assign mem_16_5_W0_clk = W0_clk;
  assign mem_16_5_W0_data = W0_data[47:40];
  assign mem_16_5_W0_en = W0_en & W0_addr_sel == 8'h10;
  assign mem_16_5_W0_mask = W0_mask[5];
  assign mem_16_6_R0_addr = R0_addr[25:0];
  assign mem_16_6_R0_clk = R0_clk;
  assign mem_16_6_R0_en = R0_en & R0_addr_sel == 8'h10;
  assign mem_16_6_W0_addr = W0_addr[25:0];
  assign mem_16_6_W0_clk = W0_clk;
  assign mem_16_6_W0_data = W0_data[55:48];
  assign mem_16_6_W0_en = W0_en & W0_addr_sel == 8'h10;
  assign mem_16_6_W0_mask = W0_mask[6];
  assign mem_16_7_R0_addr = R0_addr[25:0];
  assign mem_16_7_R0_clk = R0_clk;
  assign mem_16_7_R0_en = R0_en & R0_addr_sel == 8'h10;
  assign mem_16_7_W0_addr = W0_addr[25:0];
  assign mem_16_7_W0_clk = W0_clk;
  assign mem_16_7_W0_data = W0_data[63:56];
  assign mem_16_7_W0_en = W0_en & W0_addr_sel == 8'h10;
  assign mem_16_7_W0_mask = W0_mask[7];
  assign mem_17_0_R0_addr = R0_addr[25:0];
  assign mem_17_0_R0_clk = R0_clk;
  assign mem_17_0_R0_en = R0_en & R0_addr_sel == 8'h11;
  assign mem_17_0_W0_addr = W0_addr[25:0];
  assign mem_17_0_W0_clk = W0_clk;
  assign mem_17_0_W0_data = W0_data[7:0];
  assign mem_17_0_W0_en = W0_en & W0_addr_sel == 8'h11;
  assign mem_17_0_W0_mask = W0_mask[0];
  assign mem_17_1_R0_addr = R0_addr[25:0];
  assign mem_17_1_R0_clk = R0_clk;
  assign mem_17_1_R0_en = R0_en & R0_addr_sel == 8'h11;
  assign mem_17_1_W0_addr = W0_addr[25:0];
  assign mem_17_1_W0_clk = W0_clk;
  assign mem_17_1_W0_data = W0_data[15:8];
  assign mem_17_1_W0_en = W0_en & W0_addr_sel == 8'h11;
  assign mem_17_1_W0_mask = W0_mask[1];
  assign mem_17_2_R0_addr = R0_addr[25:0];
  assign mem_17_2_R0_clk = R0_clk;
  assign mem_17_2_R0_en = R0_en & R0_addr_sel == 8'h11;
  assign mem_17_2_W0_addr = W0_addr[25:0];
  assign mem_17_2_W0_clk = W0_clk;
  assign mem_17_2_W0_data = W0_data[23:16];
  assign mem_17_2_W0_en = W0_en & W0_addr_sel == 8'h11;
  assign mem_17_2_W0_mask = W0_mask[2];
  assign mem_17_3_R0_addr = R0_addr[25:0];
  assign mem_17_3_R0_clk = R0_clk;
  assign mem_17_3_R0_en = R0_en & R0_addr_sel == 8'h11;
  assign mem_17_3_W0_addr = W0_addr[25:0];
  assign mem_17_3_W0_clk = W0_clk;
  assign mem_17_3_W0_data = W0_data[31:24];
  assign mem_17_3_W0_en = W0_en & W0_addr_sel == 8'h11;
  assign mem_17_3_W0_mask = W0_mask[3];
  assign mem_17_4_R0_addr = R0_addr[25:0];
  assign mem_17_4_R0_clk = R0_clk;
  assign mem_17_4_R0_en = R0_en & R0_addr_sel == 8'h11;
  assign mem_17_4_W0_addr = W0_addr[25:0];
  assign mem_17_4_W0_clk = W0_clk;
  assign mem_17_4_W0_data = W0_data[39:32];
  assign mem_17_4_W0_en = W0_en & W0_addr_sel == 8'h11;
  assign mem_17_4_W0_mask = W0_mask[4];
  assign mem_17_5_R0_addr = R0_addr[25:0];
  assign mem_17_5_R0_clk = R0_clk;
  assign mem_17_5_R0_en = R0_en & R0_addr_sel == 8'h11;
  assign mem_17_5_W0_addr = W0_addr[25:0];
  assign mem_17_5_W0_clk = W0_clk;
  assign mem_17_5_W0_data = W0_data[47:40];
  assign mem_17_5_W0_en = W0_en & W0_addr_sel == 8'h11;
  assign mem_17_5_W0_mask = W0_mask[5];
  assign mem_17_6_R0_addr = R0_addr[25:0];
  assign mem_17_6_R0_clk = R0_clk;
  assign mem_17_6_R0_en = R0_en & R0_addr_sel == 8'h11;
  assign mem_17_6_W0_addr = W0_addr[25:0];
  assign mem_17_6_W0_clk = W0_clk;
  assign mem_17_6_W0_data = W0_data[55:48];
  assign mem_17_6_W0_en = W0_en & W0_addr_sel == 8'h11;
  assign mem_17_6_W0_mask = W0_mask[6];
  assign mem_17_7_R0_addr = R0_addr[25:0];
  assign mem_17_7_R0_clk = R0_clk;
  assign mem_17_7_R0_en = R0_en & R0_addr_sel == 8'h11;
  assign mem_17_7_W0_addr = W0_addr[25:0];
  assign mem_17_7_W0_clk = W0_clk;
  assign mem_17_7_W0_data = W0_data[63:56];
  assign mem_17_7_W0_en = W0_en & W0_addr_sel == 8'h11;
  assign mem_17_7_W0_mask = W0_mask[7];
  assign mem_18_0_R0_addr = R0_addr[25:0];
  assign mem_18_0_R0_clk = R0_clk;
  assign mem_18_0_R0_en = R0_en & R0_addr_sel == 8'h12;
  assign mem_18_0_W0_addr = W0_addr[25:0];
  assign mem_18_0_W0_clk = W0_clk;
  assign mem_18_0_W0_data = W0_data[7:0];
  assign mem_18_0_W0_en = W0_en & W0_addr_sel == 8'h12;
  assign mem_18_0_W0_mask = W0_mask[0];
  assign mem_18_1_R0_addr = R0_addr[25:0];
  assign mem_18_1_R0_clk = R0_clk;
  assign mem_18_1_R0_en = R0_en & R0_addr_sel == 8'h12;
  assign mem_18_1_W0_addr = W0_addr[25:0];
  assign mem_18_1_W0_clk = W0_clk;
  assign mem_18_1_W0_data = W0_data[15:8];
  assign mem_18_1_W0_en = W0_en & W0_addr_sel == 8'h12;
  assign mem_18_1_W0_mask = W0_mask[1];
  assign mem_18_2_R0_addr = R0_addr[25:0];
  assign mem_18_2_R0_clk = R0_clk;
  assign mem_18_2_R0_en = R0_en & R0_addr_sel == 8'h12;
  assign mem_18_2_W0_addr = W0_addr[25:0];
  assign mem_18_2_W0_clk = W0_clk;
  assign mem_18_2_W0_data = W0_data[23:16];
  assign mem_18_2_W0_en = W0_en & W0_addr_sel == 8'h12;
  assign mem_18_2_W0_mask = W0_mask[2];
  assign mem_18_3_R0_addr = R0_addr[25:0];
  assign mem_18_3_R0_clk = R0_clk;
  assign mem_18_3_R0_en = R0_en & R0_addr_sel == 8'h12;
  assign mem_18_3_W0_addr = W0_addr[25:0];
  assign mem_18_3_W0_clk = W0_clk;
  assign mem_18_3_W0_data = W0_data[31:24];
  assign mem_18_3_W0_en = W0_en & W0_addr_sel == 8'h12;
  assign mem_18_3_W0_mask = W0_mask[3];
  assign mem_18_4_R0_addr = R0_addr[25:0];
  assign mem_18_4_R0_clk = R0_clk;
  assign mem_18_4_R0_en = R0_en & R0_addr_sel == 8'h12;
  assign mem_18_4_W0_addr = W0_addr[25:0];
  assign mem_18_4_W0_clk = W0_clk;
  assign mem_18_4_W0_data = W0_data[39:32];
  assign mem_18_4_W0_en = W0_en & W0_addr_sel == 8'h12;
  assign mem_18_4_W0_mask = W0_mask[4];
  assign mem_18_5_R0_addr = R0_addr[25:0];
  assign mem_18_5_R0_clk = R0_clk;
  assign mem_18_5_R0_en = R0_en & R0_addr_sel == 8'h12;
  assign mem_18_5_W0_addr = W0_addr[25:0];
  assign mem_18_5_W0_clk = W0_clk;
  assign mem_18_5_W0_data = W0_data[47:40];
  assign mem_18_5_W0_en = W0_en & W0_addr_sel == 8'h12;
  assign mem_18_5_W0_mask = W0_mask[5];
  assign mem_18_6_R0_addr = R0_addr[25:0];
  assign mem_18_6_R0_clk = R0_clk;
  assign mem_18_6_R0_en = R0_en & R0_addr_sel == 8'h12;
  assign mem_18_6_W0_addr = W0_addr[25:0];
  assign mem_18_6_W0_clk = W0_clk;
  assign mem_18_6_W0_data = W0_data[55:48];
  assign mem_18_6_W0_en = W0_en & W0_addr_sel == 8'h12;
  assign mem_18_6_W0_mask = W0_mask[6];
  assign mem_18_7_R0_addr = R0_addr[25:0];
  assign mem_18_7_R0_clk = R0_clk;
  assign mem_18_7_R0_en = R0_en & R0_addr_sel == 8'h12;
  assign mem_18_7_W0_addr = W0_addr[25:0];
  assign mem_18_7_W0_clk = W0_clk;
  assign mem_18_7_W0_data = W0_data[63:56];
  assign mem_18_7_W0_en = W0_en & W0_addr_sel == 8'h12;
  assign mem_18_7_W0_mask = W0_mask[7];
  assign mem_19_0_R0_addr = R0_addr[25:0];
  assign mem_19_0_R0_clk = R0_clk;
  assign mem_19_0_R0_en = R0_en & R0_addr_sel == 8'h13;
  assign mem_19_0_W0_addr = W0_addr[25:0];
  assign mem_19_0_W0_clk = W0_clk;
  assign mem_19_0_W0_data = W0_data[7:0];
  assign mem_19_0_W0_en = W0_en & W0_addr_sel == 8'h13;
  assign mem_19_0_W0_mask = W0_mask[0];
  assign mem_19_1_R0_addr = R0_addr[25:0];
  assign mem_19_1_R0_clk = R0_clk;
  assign mem_19_1_R0_en = R0_en & R0_addr_sel == 8'h13;
  assign mem_19_1_W0_addr = W0_addr[25:0];
  assign mem_19_1_W0_clk = W0_clk;
  assign mem_19_1_W0_data = W0_data[15:8];
  assign mem_19_1_W0_en = W0_en & W0_addr_sel == 8'h13;
  assign mem_19_1_W0_mask = W0_mask[1];
  assign mem_19_2_R0_addr = R0_addr[25:0];
  assign mem_19_2_R0_clk = R0_clk;
  assign mem_19_2_R0_en = R0_en & R0_addr_sel == 8'h13;
  assign mem_19_2_W0_addr = W0_addr[25:0];
  assign mem_19_2_W0_clk = W0_clk;
  assign mem_19_2_W0_data = W0_data[23:16];
  assign mem_19_2_W0_en = W0_en & W0_addr_sel == 8'h13;
  assign mem_19_2_W0_mask = W0_mask[2];
  assign mem_19_3_R0_addr = R0_addr[25:0];
  assign mem_19_3_R0_clk = R0_clk;
  assign mem_19_3_R0_en = R0_en & R0_addr_sel == 8'h13;
  assign mem_19_3_W0_addr = W0_addr[25:0];
  assign mem_19_3_W0_clk = W0_clk;
  assign mem_19_3_W0_data = W0_data[31:24];
  assign mem_19_3_W0_en = W0_en & W0_addr_sel == 8'h13;
  assign mem_19_3_W0_mask = W0_mask[3];
  assign mem_19_4_R0_addr = R0_addr[25:0];
  assign mem_19_4_R0_clk = R0_clk;
  assign mem_19_4_R0_en = R0_en & R0_addr_sel == 8'h13;
  assign mem_19_4_W0_addr = W0_addr[25:0];
  assign mem_19_4_W0_clk = W0_clk;
  assign mem_19_4_W0_data = W0_data[39:32];
  assign mem_19_4_W0_en = W0_en & W0_addr_sel == 8'h13;
  assign mem_19_4_W0_mask = W0_mask[4];
  assign mem_19_5_R0_addr = R0_addr[25:0];
  assign mem_19_5_R0_clk = R0_clk;
  assign mem_19_5_R0_en = R0_en & R0_addr_sel == 8'h13;
  assign mem_19_5_W0_addr = W0_addr[25:0];
  assign mem_19_5_W0_clk = W0_clk;
  assign mem_19_5_W0_data = W0_data[47:40];
  assign mem_19_5_W0_en = W0_en & W0_addr_sel == 8'h13;
  assign mem_19_5_W0_mask = W0_mask[5];
  assign mem_19_6_R0_addr = R0_addr[25:0];
  assign mem_19_6_R0_clk = R0_clk;
  assign mem_19_6_R0_en = R0_en & R0_addr_sel == 8'h13;
  assign mem_19_6_W0_addr = W0_addr[25:0];
  assign mem_19_6_W0_clk = W0_clk;
  assign mem_19_6_W0_data = W0_data[55:48];
  assign mem_19_6_W0_en = W0_en & W0_addr_sel == 8'h13;
  assign mem_19_6_W0_mask = W0_mask[6];
  assign mem_19_7_R0_addr = R0_addr[25:0];
  assign mem_19_7_R0_clk = R0_clk;
  assign mem_19_7_R0_en = R0_en & R0_addr_sel == 8'h13;
  assign mem_19_7_W0_addr = W0_addr[25:0];
  assign mem_19_7_W0_clk = W0_clk;
  assign mem_19_7_W0_data = W0_data[63:56];
  assign mem_19_7_W0_en = W0_en & W0_addr_sel == 8'h13;
  assign mem_19_7_W0_mask = W0_mask[7];
  assign mem_20_0_R0_addr = R0_addr[25:0];
  assign mem_20_0_R0_clk = R0_clk;
  assign mem_20_0_R0_en = R0_en & R0_addr_sel == 8'h14;
  assign mem_20_0_W0_addr = W0_addr[25:0];
  assign mem_20_0_W0_clk = W0_clk;
  assign mem_20_0_W0_data = W0_data[7:0];
  assign mem_20_0_W0_en = W0_en & W0_addr_sel == 8'h14;
  assign mem_20_0_W0_mask = W0_mask[0];
  assign mem_20_1_R0_addr = R0_addr[25:0];
  assign mem_20_1_R0_clk = R0_clk;
  assign mem_20_1_R0_en = R0_en & R0_addr_sel == 8'h14;
  assign mem_20_1_W0_addr = W0_addr[25:0];
  assign mem_20_1_W0_clk = W0_clk;
  assign mem_20_1_W0_data = W0_data[15:8];
  assign mem_20_1_W0_en = W0_en & W0_addr_sel == 8'h14;
  assign mem_20_1_W0_mask = W0_mask[1];
  assign mem_20_2_R0_addr = R0_addr[25:0];
  assign mem_20_2_R0_clk = R0_clk;
  assign mem_20_2_R0_en = R0_en & R0_addr_sel == 8'h14;
  assign mem_20_2_W0_addr = W0_addr[25:0];
  assign mem_20_2_W0_clk = W0_clk;
  assign mem_20_2_W0_data = W0_data[23:16];
  assign mem_20_2_W0_en = W0_en & W0_addr_sel == 8'h14;
  assign mem_20_2_W0_mask = W0_mask[2];
  assign mem_20_3_R0_addr = R0_addr[25:0];
  assign mem_20_3_R0_clk = R0_clk;
  assign mem_20_3_R0_en = R0_en & R0_addr_sel == 8'h14;
  assign mem_20_3_W0_addr = W0_addr[25:0];
  assign mem_20_3_W0_clk = W0_clk;
  assign mem_20_3_W0_data = W0_data[31:24];
  assign mem_20_3_W0_en = W0_en & W0_addr_sel == 8'h14;
  assign mem_20_3_W0_mask = W0_mask[3];
  assign mem_20_4_R0_addr = R0_addr[25:0];
  assign mem_20_4_R0_clk = R0_clk;
  assign mem_20_4_R0_en = R0_en & R0_addr_sel == 8'h14;
  assign mem_20_4_W0_addr = W0_addr[25:0];
  assign mem_20_4_W0_clk = W0_clk;
  assign mem_20_4_W0_data = W0_data[39:32];
  assign mem_20_4_W0_en = W0_en & W0_addr_sel == 8'h14;
  assign mem_20_4_W0_mask = W0_mask[4];
  assign mem_20_5_R0_addr = R0_addr[25:0];
  assign mem_20_5_R0_clk = R0_clk;
  assign mem_20_5_R0_en = R0_en & R0_addr_sel == 8'h14;
  assign mem_20_5_W0_addr = W0_addr[25:0];
  assign mem_20_5_W0_clk = W0_clk;
  assign mem_20_5_W0_data = W0_data[47:40];
  assign mem_20_5_W0_en = W0_en & W0_addr_sel == 8'h14;
  assign mem_20_5_W0_mask = W0_mask[5];
  assign mem_20_6_R0_addr = R0_addr[25:0];
  assign mem_20_6_R0_clk = R0_clk;
  assign mem_20_6_R0_en = R0_en & R0_addr_sel == 8'h14;
  assign mem_20_6_W0_addr = W0_addr[25:0];
  assign mem_20_6_W0_clk = W0_clk;
  assign mem_20_6_W0_data = W0_data[55:48];
  assign mem_20_6_W0_en = W0_en & W0_addr_sel == 8'h14;
  assign mem_20_6_W0_mask = W0_mask[6];
  assign mem_20_7_R0_addr = R0_addr[25:0];
  assign mem_20_7_R0_clk = R0_clk;
  assign mem_20_7_R0_en = R0_en & R0_addr_sel == 8'h14;
  assign mem_20_7_W0_addr = W0_addr[25:0];
  assign mem_20_7_W0_clk = W0_clk;
  assign mem_20_7_W0_data = W0_data[63:56];
  assign mem_20_7_W0_en = W0_en & W0_addr_sel == 8'h14;
  assign mem_20_7_W0_mask = W0_mask[7];
  assign mem_21_0_R0_addr = R0_addr[25:0];
  assign mem_21_0_R0_clk = R0_clk;
  assign mem_21_0_R0_en = R0_en & R0_addr_sel == 8'h15;
  assign mem_21_0_W0_addr = W0_addr[25:0];
  assign mem_21_0_W0_clk = W0_clk;
  assign mem_21_0_W0_data = W0_data[7:0];
  assign mem_21_0_W0_en = W0_en & W0_addr_sel == 8'h15;
  assign mem_21_0_W0_mask = W0_mask[0];
  assign mem_21_1_R0_addr = R0_addr[25:0];
  assign mem_21_1_R0_clk = R0_clk;
  assign mem_21_1_R0_en = R0_en & R0_addr_sel == 8'h15;
  assign mem_21_1_W0_addr = W0_addr[25:0];
  assign mem_21_1_W0_clk = W0_clk;
  assign mem_21_1_W0_data = W0_data[15:8];
  assign mem_21_1_W0_en = W0_en & W0_addr_sel == 8'h15;
  assign mem_21_1_W0_mask = W0_mask[1];
  assign mem_21_2_R0_addr = R0_addr[25:0];
  assign mem_21_2_R0_clk = R0_clk;
  assign mem_21_2_R0_en = R0_en & R0_addr_sel == 8'h15;
  assign mem_21_2_W0_addr = W0_addr[25:0];
  assign mem_21_2_W0_clk = W0_clk;
  assign mem_21_2_W0_data = W0_data[23:16];
  assign mem_21_2_W0_en = W0_en & W0_addr_sel == 8'h15;
  assign mem_21_2_W0_mask = W0_mask[2];
  assign mem_21_3_R0_addr = R0_addr[25:0];
  assign mem_21_3_R0_clk = R0_clk;
  assign mem_21_3_R0_en = R0_en & R0_addr_sel == 8'h15;
  assign mem_21_3_W0_addr = W0_addr[25:0];
  assign mem_21_3_W0_clk = W0_clk;
  assign mem_21_3_W0_data = W0_data[31:24];
  assign mem_21_3_W0_en = W0_en & W0_addr_sel == 8'h15;
  assign mem_21_3_W0_mask = W0_mask[3];
  assign mem_21_4_R0_addr = R0_addr[25:0];
  assign mem_21_4_R0_clk = R0_clk;
  assign mem_21_4_R0_en = R0_en & R0_addr_sel == 8'h15;
  assign mem_21_4_W0_addr = W0_addr[25:0];
  assign mem_21_4_W0_clk = W0_clk;
  assign mem_21_4_W0_data = W0_data[39:32];
  assign mem_21_4_W0_en = W0_en & W0_addr_sel == 8'h15;
  assign mem_21_4_W0_mask = W0_mask[4];
  assign mem_21_5_R0_addr = R0_addr[25:0];
  assign mem_21_5_R0_clk = R0_clk;
  assign mem_21_5_R0_en = R0_en & R0_addr_sel == 8'h15;
  assign mem_21_5_W0_addr = W0_addr[25:0];
  assign mem_21_5_W0_clk = W0_clk;
  assign mem_21_5_W0_data = W0_data[47:40];
  assign mem_21_5_W0_en = W0_en & W0_addr_sel == 8'h15;
  assign mem_21_5_W0_mask = W0_mask[5];
  assign mem_21_6_R0_addr = R0_addr[25:0];
  assign mem_21_6_R0_clk = R0_clk;
  assign mem_21_6_R0_en = R0_en & R0_addr_sel == 8'h15;
  assign mem_21_6_W0_addr = W0_addr[25:0];
  assign mem_21_6_W0_clk = W0_clk;
  assign mem_21_6_W0_data = W0_data[55:48];
  assign mem_21_6_W0_en = W0_en & W0_addr_sel == 8'h15;
  assign mem_21_6_W0_mask = W0_mask[6];
  assign mem_21_7_R0_addr = R0_addr[25:0];
  assign mem_21_7_R0_clk = R0_clk;
  assign mem_21_7_R0_en = R0_en & R0_addr_sel == 8'h15;
  assign mem_21_7_W0_addr = W0_addr[25:0];
  assign mem_21_7_W0_clk = W0_clk;
  assign mem_21_7_W0_data = W0_data[63:56];
  assign mem_21_7_W0_en = W0_en & W0_addr_sel == 8'h15;
  assign mem_21_7_W0_mask = W0_mask[7];
  assign mem_22_0_R0_addr = R0_addr[25:0];
  assign mem_22_0_R0_clk = R0_clk;
  assign mem_22_0_R0_en = R0_en & R0_addr_sel == 8'h16;
  assign mem_22_0_W0_addr = W0_addr[25:0];
  assign mem_22_0_W0_clk = W0_clk;
  assign mem_22_0_W0_data = W0_data[7:0];
  assign mem_22_0_W0_en = W0_en & W0_addr_sel == 8'h16;
  assign mem_22_0_W0_mask = W0_mask[0];
  assign mem_22_1_R0_addr = R0_addr[25:0];
  assign mem_22_1_R0_clk = R0_clk;
  assign mem_22_1_R0_en = R0_en & R0_addr_sel == 8'h16;
  assign mem_22_1_W0_addr = W0_addr[25:0];
  assign mem_22_1_W0_clk = W0_clk;
  assign mem_22_1_W0_data = W0_data[15:8];
  assign mem_22_1_W0_en = W0_en & W0_addr_sel == 8'h16;
  assign mem_22_1_W0_mask = W0_mask[1];
  assign mem_22_2_R0_addr = R0_addr[25:0];
  assign mem_22_2_R0_clk = R0_clk;
  assign mem_22_2_R0_en = R0_en & R0_addr_sel == 8'h16;
  assign mem_22_2_W0_addr = W0_addr[25:0];
  assign mem_22_2_W0_clk = W0_clk;
  assign mem_22_2_W0_data = W0_data[23:16];
  assign mem_22_2_W0_en = W0_en & W0_addr_sel == 8'h16;
  assign mem_22_2_W0_mask = W0_mask[2];
  assign mem_22_3_R0_addr = R0_addr[25:0];
  assign mem_22_3_R0_clk = R0_clk;
  assign mem_22_3_R0_en = R0_en & R0_addr_sel == 8'h16;
  assign mem_22_3_W0_addr = W0_addr[25:0];
  assign mem_22_3_W0_clk = W0_clk;
  assign mem_22_3_W0_data = W0_data[31:24];
  assign mem_22_3_W0_en = W0_en & W0_addr_sel == 8'h16;
  assign mem_22_3_W0_mask = W0_mask[3];
  assign mem_22_4_R0_addr = R0_addr[25:0];
  assign mem_22_4_R0_clk = R0_clk;
  assign mem_22_4_R0_en = R0_en & R0_addr_sel == 8'h16;
  assign mem_22_4_W0_addr = W0_addr[25:0];
  assign mem_22_4_W0_clk = W0_clk;
  assign mem_22_4_W0_data = W0_data[39:32];
  assign mem_22_4_W0_en = W0_en & W0_addr_sel == 8'h16;
  assign mem_22_4_W0_mask = W0_mask[4];
  assign mem_22_5_R0_addr = R0_addr[25:0];
  assign mem_22_5_R0_clk = R0_clk;
  assign mem_22_5_R0_en = R0_en & R0_addr_sel == 8'h16;
  assign mem_22_5_W0_addr = W0_addr[25:0];
  assign mem_22_5_W0_clk = W0_clk;
  assign mem_22_5_W0_data = W0_data[47:40];
  assign mem_22_5_W0_en = W0_en & W0_addr_sel == 8'h16;
  assign mem_22_5_W0_mask = W0_mask[5];
  assign mem_22_6_R0_addr = R0_addr[25:0];
  assign mem_22_6_R0_clk = R0_clk;
  assign mem_22_6_R0_en = R0_en & R0_addr_sel == 8'h16;
  assign mem_22_6_W0_addr = W0_addr[25:0];
  assign mem_22_6_W0_clk = W0_clk;
  assign mem_22_6_W0_data = W0_data[55:48];
  assign mem_22_6_W0_en = W0_en & W0_addr_sel == 8'h16;
  assign mem_22_6_W0_mask = W0_mask[6];
  assign mem_22_7_R0_addr = R0_addr[25:0];
  assign mem_22_7_R0_clk = R0_clk;
  assign mem_22_7_R0_en = R0_en & R0_addr_sel == 8'h16;
  assign mem_22_7_W0_addr = W0_addr[25:0];
  assign mem_22_7_W0_clk = W0_clk;
  assign mem_22_7_W0_data = W0_data[63:56];
  assign mem_22_7_W0_en = W0_en & W0_addr_sel == 8'h16;
  assign mem_22_7_W0_mask = W0_mask[7];
  assign mem_23_0_R0_addr = R0_addr[25:0];
  assign mem_23_0_R0_clk = R0_clk;
  assign mem_23_0_R0_en = R0_en & R0_addr_sel == 8'h17;
  assign mem_23_0_W0_addr = W0_addr[25:0];
  assign mem_23_0_W0_clk = W0_clk;
  assign mem_23_0_W0_data = W0_data[7:0];
  assign mem_23_0_W0_en = W0_en & W0_addr_sel == 8'h17;
  assign mem_23_0_W0_mask = W0_mask[0];
  assign mem_23_1_R0_addr = R0_addr[25:0];
  assign mem_23_1_R0_clk = R0_clk;
  assign mem_23_1_R0_en = R0_en & R0_addr_sel == 8'h17;
  assign mem_23_1_W0_addr = W0_addr[25:0];
  assign mem_23_1_W0_clk = W0_clk;
  assign mem_23_1_W0_data = W0_data[15:8];
  assign mem_23_1_W0_en = W0_en & W0_addr_sel == 8'h17;
  assign mem_23_1_W0_mask = W0_mask[1];
  assign mem_23_2_R0_addr = R0_addr[25:0];
  assign mem_23_2_R0_clk = R0_clk;
  assign mem_23_2_R0_en = R0_en & R0_addr_sel == 8'h17;
  assign mem_23_2_W0_addr = W0_addr[25:0];
  assign mem_23_2_W0_clk = W0_clk;
  assign mem_23_2_W0_data = W0_data[23:16];
  assign mem_23_2_W0_en = W0_en & W0_addr_sel == 8'h17;
  assign mem_23_2_W0_mask = W0_mask[2];
  assign mem_23_3_R0_addr = R0_addr[25:0];
  assign mem_23_3_R0_clk = R0_clk;
  assign mem_23_3_R0_en = R0_en & R0_addr_sel == 8'h17;
  assign mem_23_3_W0_addr = W0_addr[25:0];
  assign mem_23_3_W0_clk = W0_clk;
  assign mem_23_3_W0_data = W0_data[31:24];
  assign mem_23_3_W0_en = W0_en & W0_addr_sel == 8'h17;
  assign mem_23_3_W0_mask = W0_mask[3];
  assign mem_23_4_R0_addr = R0_addr[25:0];
  assign mem_23_4_R0_clk = R0_clk;
  assign mem_23_4_R0_en = R0_en & R0_addr_sel == 8'h17;
  assign mem_23_4_W0_addr = W0_addr[25:0];
  assign mem_23_4_W0_clk = W0_clk;
  assign mem_23_4_W0_data = W0_data[39:32];
  assign mem_23_4_W0_en = W0_en & W0_addr_sel == 8'h17;
  assign mem_23_4_W0_mask = W0_mask[4];
  assign mem_23_5_R0_addr = R0_addr[25:0];
  assign mem_23_5_R0_clk = R0_clk;
  assign mem_23_5_R0_en = R0_en & R0_addr_sel == 8'h17;
  assign mem_23_5_W0_addr = W0_addr[25:0];
  assign mem_23_5_W0_clk = W0_clk;
  assign mem_23_5_W0_data = W0_data[47:40];
  assign mem_23_5_W0_en = W0_en & W0_addr_sel == 8'h17;
  assign mem_23_5_W0_mask = W0_mask[5];
  assign mem_23_6_R0_addr = R0_addr[25:0];
  assign mem_23_6_R0_clk = R0_clk;
  assign mem_23_6_R0_en = R0_en & R0_addr_sel == 8'h17;
  assign mem_23_6_W0_addr = W0_addr[25:0];
  assign mem_23_6_W0_clk = W0_clk;
  assign mem_23_6_W0_data = W0_data[55:48];
  assign mem_23_6_W0_en = W0_en & W0_addr_sel == 8'h17;
  assign mem_23_6_W0_mask = W0_mask[6];
  assign mem_23_7_R0_addr = R0_addr[25:0];
  assign mem_23_7_R0_clk = R0_clk;
  assign mem_23_7_R0_en = R0_en & R0_addr_sel == 8'h17;
  assign mem_23_7_W0_addr = W0_addr[25:0];
  assign mem_23_7_W0_clk = W0_clk;
  assign mem_23_7_W0_data = W0_data[63:56];
  assign mem_23_7_W0_en = W0_en & W0_addr_sel == 8'h17;
  assign mem_23_7_W0_mask = W0_mask[7];
  assign mem_24_0_R0_addr = R0_addr[25:0];
  assign mem_24_0_R0_clk = R0_clk;
  assign mem_24_0_R0_en = R0_en & R0_addr_sel == 8'h18;
  assign mem_24_0_W0_addr = W0_addr[25:0];
  assign mem_24_0_W0_clk = W0_clk;
  assign mem_24_0_W0_data = W0_data[7:0];
  assign mem_24_0_W0_en = W0_en & W0_addr_sel == 8'h18;
  assign mem_24_0_W0_mask = W0_mask[0];
  assign mem_24_1_R0_addr = R0_addr[25:0];
  assign mem_24_1_R0_clk = R0_clk;
  assign mem_24_1_R0_en = R0_en & R0_addr_sel == 8'h18;
  assign mem_24_1_W0_addr = W0_addr[25:0];
  assign mem_24_1_W0_clk = W0_clk;
  assign mem_24_1_W0_data = W0_data[15:8];
  assign mem_24_1_W0_en = W0_en & W0_addr_sel == 8'h18;
  assign mem_24_1_W0_mask = W0_mask[1];
  assign mem_24_2_R0_addr = R0_addr[25:0];
  assign mem_24_2_R0_clk = R0_clk;
  assign mem_24_2_R0_en = R0_en & R0_addr_sel == 8'h18;
  assign mem_24_2_W0_addr = W0_addr[25:0];
  assign mem_24_2_W0_clk = W0_clk;
  assign mem_24_2_W0_data = W0_data[23:16];
  assign mem_24_2_W0_en = W0_en & W0_addr_sel == 8'h18;
  assign mem_24_2_W0_mask = W0_mask[2];
  assign mem_24_3_R0_addr = R0_addr[25:0];
  assign mem_24_3_R0_clk = R0_clk;
  assign mem_24_3_R0_en = R0_en & R0_addr_sel == 8'h18;
  assign mem_24_3_W0_addr = W0_addr[25:0];
  assign mem_24_3_W0_clk = W0_clk;
  assign mem_24_3_W0_data = W0_data[31:24];
  assign mem_24_3_W0_en = W0_en & W0_addr_sel == 8'h18;
  assign mem_24_3_W0_mask = W0_mask[3];
  assign mem_24_4_R0_addr = R0_addr[25:0];
  assign mem_24_4_R0_clk = R0_clk;
  assign mem_24_4_R0_en = R0_en & R0_addr_sel == 8'h18;
  assign mem_24_4_W0_addr = W0_addr[25:0];
  assign mem_24_4_W0_clk = W0_clk;
  assign mem_24_4_W0_data = W0_data[39:32];
  assign mem_24_4_W0_en = W0_en & W0_addr_sel == 8'h18;
  assign mem_24_4_W0_mask = W0_mask[4];
  assign mem_24_5_R0_addr = R0_addr[25:0];
  assign mem_24_5_R0_clk = R0_clk;
  assign mem_24_5_R0_en = R0_en & R0_addr_sel == 8'h18;
  assign mem_24_5_W0_addr = W0_addr[25:0];
  assign mem_24_5_W0_clk = W0_clk;
  assign mem_24_5_W0_data = W0_data[47:40];
  assign mem_24_5_W0_en = W0_en & W0_addr_sel == 8'h18;
  assign mem_24_5_W0_mask = W0_mask[5];
  assign mem_24_6_R0_addr = R0_addr[25:0];
  assign mem_24_6_R0_clk = R0_clk;
  assign mem_24_6_R0_en = R0_en & R0_addr_sel == 8'h18;
  assign mem_24_6_W0_addr = W0_addr[25:0];
  assign mem_24_6_W0_clk = W0_clk;
  assign mem_24_6_W0_data = W0_data[55:48];
  assign mem_24_6_W0_en = W0_en & W0_addr_sel == 8'h18;
  assign mem_24_6_W0_mask = W0_mask[6];
  assign mem_24_7_R0_addr = R0_addr[25:0];
  assign mem_24_7_R0_clk = R0_clk;
  assign mem_24_7_R0_en = R0_en & R0_addr_sel == 8'h18;
  assign mem_24_7_W0_addr = W0_addr[25:0];
  assign mem_24_7_W0_clk = W0_clk;
  assign mem_24_7_W0_data = W0_data[63:56];
  assign mem_24_7_W0_en = W0_en & W0_addr_sel == 8'h18;
  assign mem_24_7_W0_mask = W0_mask[7];
  assign mem_25_0_R0_addr = R0_addr[25:0];
  assign mem_25_0_R0_clk = R0_clk;
  assign mem_25_0_R0_en = R0_en & R0_addr_sel == 8'h19;
  assign mem_25_0_W0_addr = W0_addr[25:0];
  assign mem_25_0_W0_clk = W0_clk;
  assign mem_25_0_W0_data = W0_data[7:0];
  assign mem_25_0_W0_en = W0_en & W0_addr_sel == 8'h19;
  assign mem_25_0_W0_mask = W0_mask[0];
  assign mem_25_1_R0_addr = R0_addr[25:0];
  assign mem_25_1_R0_clk = R0_clk;
  assign mem_25_1_R0_en = R0_en & R0_addr_sel == 8'h19;
  assign mem_25_1_W0_addr = W0_addr[25:0];
  assign mem_25_1_W0_clk = W0_clk;
  assign mem_25_1_W0_data = W0_data[15:8];
  assign mem_25_1_W0_en = W0_en & W0_addr_sel == 8'h19;
  assign mem_25_1_W0_mask = W0_mask[1];
  assign mem_25_2_R0_addr = R0_addr[25:0];
  assign mem_25_2_R0_clk = R0_clk;
  assign mem_25_2_R0_en = R0_en & R0_addr_sel == 8'h19;
  assign mem_25_2_W0_addr = W0_addr[25:0];
  assign mem_25_2_W0_clk = W0_clk;
  assign mem_25_2_W0_data = W0_data[23:16];
  assign mem_25_2_W0_en = W0_en & W0_addr_sel == 8'h19;
  assign mem_25_2_W0_mask = W0_mask[2];
  assign mem_25_3_R0_addr = R0_addr[25:0];
  assign mem_25_3_R0_clk = R0_clk;
  assign mem_25_3_R0_en = R0_en & R0_addr_sel == 8'h19;
  assign mem_25_3_W0_addr = W0_addr[25:0];
  assign mem_25_3_W0_clk = W0_clk;
  assign mem_25_3_W0_data = W0_data[31:24];
  assign mem_25_3_W0_en = W0_en & W0_addr_sel == 8'h19;
  assign mem_25_3_W0_mask = W0_mask[3];
  assign mem_25_4_R0_addr = R0_addr[25:0];
  assign mem_25_4_R0_clk = R0_clk;
  assign mem_25_4_R0_en = R0_en & R0_addr_sel == 8'h19;
  assign mem_25_4_W0_addr = W0_addr[25:0];
  assign mem_25_4_W0_clk = W0_clk;
  assign mem_25_4_W0_data = W0_data[39:32];
  assign mem_25_4_W0_en = W0_en & W0_addr_sel == 8'h19;
  assign mem_25_4_W0_mask = W0_mask[4];
  assign mem_25_5_R0_addr = R0_addr[25:0];
  assign mem_25_5_R0_clk = R0_clk;
  assign mem_25_5_R0_en = R0_en & R0_addr_sel == 8'h19;
  assign mem_25_5_W0_addr = W0_addr[25:0];
  assign mem_25_5_W0_clk = W0_clk;
  assign mem_25_5_W0_data = W0_data[47:40];
  assign mem_25_5_W0_en = W0_en & W0_addr_sel == 8'h19;
  assign mem_25_5_W0_mask = W0_mask[5];
  assign mem_25_6_R0_addr = R0_addr[25:0];
  assign mem_25_6_R0_clk = R0_clk;
  assign mem_25_6_R0_en = R0_en & R0_addr_sel == 8'h19;
  assign mem_25_6_W0_addr = W0_addr[25:0];
  assign mem_25_6_W0_clk = W0_clk;
  assign mem_25_6_W0_data = W0_data[55:48];
  assign mem_25_6_W0_en = W0_en & W0_addr_sel == 8'h19;
  assign mem_25_6_W0_mask = W0_mask[6];
  assign mem_25_7_R0_addr = R0_addr[25:0];
  assign mem_25_7_R0_clk = R0_clk;
  assign mem_25_7_R0_en = R0_en & R0_addr_sel == 8'h19;
  assign mem_25_7_W0_addr = W0_addr[25:0];
  assign mem_25_7_W0_clk = W0_clk;
  assign mem_25_7_W0_data = W0_data[63:56];
  assign mem_25_7_W0_en = W0_en & W0_addr_sel == 8'h19;
  assign mem_25_7_W0_mask = W0_mask[7];
  assign mem_26_0_R0_addr = R0_addr[25:0];
  assign mem_26_0_R0_clk = R0_clk;
  assign mem_26_0_R0_en = R0_en & R0_addr_sel == 8'h1a;
  assign mem_26_0_W0_addr = W0_addr[25:0];
  assign mem_26_0_W0_clk = W0_clk;
  assign mem_26_0_W0_data = W0_data[7:0];
  assign mem_26_0_W0_en = W0_en & W0_addr_sel == 8'h1a;
  assign mem_26_0_W0_mask = W0_mask[0];
  assign mem_26_1_R0_addr = R0_addr[25:0];
  assign mem_26_1_R0_clk = R0_clk;
  assign mem_26_1_R0_en = R0_en & R0_addr_sel == 8'h1a;
  assign mem_26_1_W0_addr = W0_addr[25:0];
  assign mem_26_1_W0_clk = W0_clk;
  assign mem_26_1_W0_data = W0_data[15:8];
  assign mem_26_1_W0_en = W0_en & W0_addr_sel == 8'h1a;
  assign mem_26_1_W0_mask = W0_mask[1];
  assign mem_26_2_R0_addr = R0_addr[25:0];
  assign mem_26_2_R0_clk = R0_clk;
  assign mem_26_2_R0_en = R0_en & R0_addr_sel == 8'h1a;
  assign mem_26_2_W0_addr = W0_addr[25:0];
  assign mem_26_2_W0_clk = W0_clk;
  assign mem_26_2_W0_data = W0_data[23:16];
  assign mem_26_2_W0_en = W0_en & W0_addr_sel == 8'h1a;
  assign mem_26_2_W0_mask = W0_mask[2];
  assign mem_26_3_R0_addr = R0_addr[25:0];
  assign mem_26_3_R0_clk = R0_clk;
  assign mem_26_3_R0_en = R0_en & R0_addr_sel == 8'h1a;
  assign mem_26_3_W0_addr = W0_addr[25:0];
  assign mem_26_3_W0_clk = W0_clk;
  assign mem_26_3_W0_data = W0_data[31:24];
  assign mem_26_3_W0_en = W0_en & W0_addr_sel == 8'h1a;
  assign mem_26_3_W0_mask = W0_mask[3];
  assign mem_26_4_R0_addr = R0_addr[25:0];
  assign mem_26_4_R0_clk = R0_clk;
  assign mem_26_4_R0_en = R0_en & R0_addr_sel == 8'h1a;
  assign mem_26_4_W0_addr = W0_addr[25:0];
  assign mem_26_4_W0_clk = W0_clk;
  assign mem_26_4_W0_data = W0_data[39:32];
  assign mem_26_4_W0_en = W0_en & W0_addr_sel == 8'h1a;
  assign mem_26_4_W0_mask = W0_mask[4];
  assign mem_26_5_R0_addr = R0_addr[25:0];
  assign mem_26_5_R0_clk = R0_clk;
  assign mem_26_5_R0_en = R0_en & R0_addr_sel == 8'h1a;
  assign mem_26_5_W0_addr = W0_addr[25:0];
  assign mem_26_5_W0_clk = W0_clk;
  assign mem_26_5_W0_data = W0_data[47:40];
  assign mem_26_5_W0_en = W0_en & W0_addr_sel == 8'h1a;
  assign mem_26_5_W0_mask = W0_mask[5];
  assign mem_26_6_R0_addr = R0_addr[25:0];
  assign mem_26_6_R0_clk = R0_clk;
  assign mem_26_6_R0_en = R0_en & R0_addr_sel == 8'h1a;
  assign mem_26_6_W0_addr = W0_addr[25:0];
  assign mem_26_6_W0_clk = W0_clk;
  assign mem_26_6_W0_data = W0_data[55:48];
  assign mem_26_6_W0_en = W0_en & W0_addr_sel == 8'h1a;
  assign mem_26_6_W0_mask = W0_mask[6];
  assign mem_26_7_R0_addr = R0_addr[25:0];
  assign mem_26_7_R0_clk = R0_clk;
  assign mem_26_7_R0_en = R0_en & R0_addr_sel == 8'h1a;
  assign mem_26_7_W0_addr = W0_addr[25:0];
  assign mem_26_7_W0_clk = W0_clk;
  assign mem_26_7_W0_data = W0_data[63:56];
  assign mem_26_7_W0_en = W0_en & W0_addr_sel == 8'h1a;
  assign mem_26_7_W0_mask = W0_mask[7];
  assign mem_27_0_R0_addr = R0_addr[25:0];
  assign mem_27_0_R0_clk = R0_clk;
  assign mem_27_0_R0_en = R0_en & R0_addr_sel == 8'h1b;
  assign mem_27_0_W0_addr = W0_addr[25:0];
  assign mem_27_0_W0_clk = W0_clk;
  assign mem_27_0_W0_data = W0_data[7:0];
  assign mem_27_0_W0_en = W0_en & W0_addr_sel == 8'h1b;
  assign mem_27_0_W0_mask = W0_mask[0];
  assign mem_27_1_R0_addr = R0_addr[25:0];
  assign mem_27_1_R0_clk = R0_clk;
  assign mem_27_1_R0_en = R0_en & R0_addr_sel == 8'h1b;
  assign mem_27_1_W0_addr = W0_addr[25:0];
  assign mem_27_1_W0_clk = W0_clk;
  assign mem_27_1_W0_data = W0_data[15:8];
  assign mem_27_1_W0_en = W0_en & W0_addr_sel == 8'h1b;
  assign mem_27_1_W0_mask = W0_mask[1];
  assign mem_27_2_R0_addr = R0_addr[25:0];
  assign mem_27_2_R0_clk = R0_clk;
  assign mem_27_2_R0_en = R0_en & R0_addr_sel == 8'h1b;
  assign mem_27_2_W0_addr = W0_addr[25:0];
  assign mem_27_2_W0_clk = W0_clk;
  assign mem_27_2_W0_data = W0_data[23:16];
  assign mem_27_2_W0_en = W0_en & W0_addr_sel == 8'h1b;
  assign mem_27_2_W0_mask = W0_mask[2];
  assign mem_27_3_R0_addr = R0_addr[25:0];
  assign mem_27_3_R0_clk = R0_clk;
  assign mem_27_3_R0_en = R0_en & R0_addr_sel == 8'h1b;
  assign mem_27_3_W0_addr = W0_addr[25:0];
  assign mem_27_3_W0_clk = W0_clk;
  assign mem_27_3_W0_data = W0_data[31:24];
  assign mem_27_3_W0_en = W0_en & W0_addr_sel == 8'h1b;
  assign mem_27_3_W0_mask = W0_mask[3];
  assign mem_27_4_R0_addr = R0_addr[25:0];
  assign mem_27_4_R0_clk = R0_clk;
  assign mem_27_4_R0_en = R0_en & R0_addr_sel == 8'h1b;
  assign mem_27_4_W0_addr = W0_addr[25:0];
  assign mem_27_4_W0_clk = W0_clk;
  assign mem_27_4_W0_data = W0_data[39:32];
  assign mem_27_4_W0_en = W0_en & W0_addr_sel == 8'h1b;
  assign mem_27_4_W0_mask = W0_mask[4];
  assign mem_27_5_R0_addr = R0_addr[25:0];
  assign mem_27_5_R0_clk = R0_clk;
  assign mem_27_5_R0_en = R0_en & R0_addr_sel == 8'h1b;
  assign mem_27_5_W0_addr = W0_addr[25:0];
  assign mem_27_5_W0_clk = W0_clk;
  assign mem_27_5_W0_data = W0_data[47:40];
  assign mem_27_5_W0_en = W0_en & W0_addr_sel == 8'h1b;
  assign mem_27_5_W0_mask = W0_mask[5];
  assign mem_27_6_R0_addr = R0_addr[25:0];
  assign mem_27_6_R0_clk = R0_clk;
  assign mem_27_6_R0_en = R0_en & R0_addr_sel == 8'h1b;
  assign mem_27_6_W0_addr = W0_addr[25:0];
  assign mem_27_6_W0_clk = W0_clk;
  assign mem_27_6_W0_data = W0_data[55:48];
  assign mem_27_6_W0_en = W0_en & W0_addr_sel == 8'h1b;
  assign mem_27_6_W0_mask = W0_mask[6];
  assign mem_27_7_R0_addr = R0_addr[25:0];
  assign mem_27_7_R0_clk = R0_clk;
  assign mem_27_7_R0_en = R0_en & R0_addr_sel == 8'h1b;
  assign mem_27_7_W0_addr = W0_addr[25:0];
  assign mem_27_7_W0_clk = W0_clk;
  assign mem_27_7_W0_data = W0_data[63:56];
  assign mem_27_7_W0_en = W0_en & W0_addr_sel == 8'h1b;
  assign mem_27_7_W0_mask = W0_mask[7];
  assign mem_28_0_R0_addr = R0_addr[25:0];
  assign mem_28_0_R0_clk = R0_clk;
  assign mem_28_0_R0_en = R0_en & R0_addr_sel == 8'h1c;
  assign mem_28_0_W0_addr = W0_addr[25:0];
  assign mem_28_0_W0_clk = W0_clk;
  assign mem_28_0_W0_data = W0_data[7:0];
  assign mem_28_0_W0_en = W0_en & W0_addr_sel == 8'h1c;
  assign mem_28_0_W0_mask = W0_mask[0];
  assign mem_28_1_R0_addr = R0_addr[25:0];
  assign mem_28_1_R0_clk = R0_clk;
  assign mem_28_1_R0_en = R0_en & R0_addr_sel == 8'h1c;
  assign mem_28_1_W0_addr = W0_addr[25:0];
  assign mem_28_1_W0_clk = W0_clk;
  assign mem_28_1_W0_data = W0_data[15:8];
  assign mem_28_1_W0_en = W0_en & W0_addr_sel == 8'h1c;
  assign mem_28_1_W0_mask = W0_mask[1];
  assign mem_28_2_R0_addr = R0_addr[25:0];
  assign mem_28_2_R0_clk = R0_clk;
  assign mem_28_2_R0_en = R0_en & R0_addr_sel == 8'h1c;
  assign mem_28_2_W0_addr = W0_addr[25:0];
  assign mem_28_2_W0_clk = W0_clk;
  assign mem_28_2_W0_data = W0_data[23:16];
  assign mem_28_2_W0_en = W0_en & W0_addr_sel == 8'h1c;
  assign mem_28_2_W0_mask = W0_mask[2];
  assign mem_28_3_R0_addr = R0_addr[25:0];
  assign mem_28_3_R0_clk = R0_clk;
  assign mem_28_3_R0_en = R0_en & R0_addr_sel == 8'h1c;
  assign mem_28_3_W0_addr = W0_addr[25:0];
  assign mem_28_3_W0_clk = W0_clk;
  assign mem_28_3_W0_data = W0_data[31:24];
  assign mem_28_3_W0_en = W0_en & W0_addr_sel == 8'h1c;
  assign mem_28_3_W0_mask = W0_mask[3];
  assign mem_28_4_R0_addr = R0_addr[25:0];
  assign mem_28_4_R0_clk = R0_clk;
  assign mem_28_4_R0_en = R0_en & R0_addr_sel == 8'h1c;
  assign mem_28_4_W0_addr = W0_addr[25:0];
  assign mem_28_4_W0_clk = W0_clk;
  assign mem_28_4_W0_data = W0_data[39:32];
  assign mem_28_4_W0_en = W0_en & W0_addr_sel == 8'h1c;
  assign mem_28_4_W0_mask = W0_mask[4];
  assign mem_28_5_R0_addr = R0_addr[25:0];
  assign mem_28_5_R0_clk = R0_clk;
  assign mem_28_5_R0_en = R0_en & R0_addr_sel == 8'h1c;
  assign mem_28_5_W0_addr = W0_addr[25:0];
  assign mem_28_5_W0_clk = W0_clk;
  assign mem_28_5_W0_data = W0_data[47:40];
  assign mem_28_5_W0_en = W0_en & W0_addr_sel == 8'h1c;
  assign mem_28_5_W0_mask = W0_mask[5];
  assign mem_28_6_R0_addr = R0_addr[25:0];
  assign mem_28_6_R0_clk = R0_clk;
  assign mem_28_6_R0_en = R0_en & R0_addr_sel == 8'h1c;
  assign mem_28_6_W0_addr = W0_addr[25:0];
  assign mem_28_6_W0_clk = W0_clk;
  assign mem_28_6_W0_data = W0_data[55:48];
  assign mem_28_6_W0_en = W0_en & W0_addr_sel == 8'h1c;
  assign mem_28_6_W0_mask = W0_mask[6];
  assign mem_28_7_R0_addr = R0_addr[25:0];
  assign mem_28_7_R0_clk = R0_clk;
  assign mem_28_7_R0_en = R0_en & R0_addr_sel == 8'h1c;
  assign mem_28_7_W0_addr = W0_addr[25:0];
  assign mem_28_7_W0_clk = W0_clk;
  assign mem_28_7_W0_data = W0_data[63:56];
  assign mem_28_7_W0_en = W0_en & W0_addr_sel == 8'h1c;
  assign mem_28_7_W0_mask = W0_mask[7];
  assign mem_29_0_R0_addr = R0_addr[25:0];
  assign mem_29_0_R0_clk = R0_clk;
  assign mem_29_0_R0_en = R0_en & R0_addr_sel == 8'h1d;
  assign mem_29_0_W0_addr = W0_addr[25:0];
  assign mem_29_0_W0_clk = W0_clk;
  assign mem_29_0_W0_data = W0_data[7:0];
  assign mem_29_0_W0_en = W0_en & W0_addr_sel == 8'h1d;
  assign mem_29_0_W0_mask = W0_mask[0];
  assign mem_29_1_R0_addr = R0_addr[25:0];
  assign mem_29_1_R0_clk = R0_clk;
  assign mem_29_1_R0_en = R0_en & R0_addr_sel == 8'h1d;
  assign mem_29_1_W0_addr = W0_addr[25:0];
  assign mem_29_1_W0_clk = W0_clk;
  assign mem_29_1_W0_data = W0_data[15:8];
  assign mem_29_1_W0_en = W0_en & W0_addr_sel == 8'h1d;
  assign mem_29_1_W0_mask = W0_mask[1];
  assign mem_29_2_R0_addr = R0_addr[25:0];
  assign mem_29_2_R0_clk = R0_clk;
  assign mem_29_2_R0_en = R0_en & R0_addr_sel == 8'h1d;
  assign mem_29_2_W0_addr = W0_addr[25:0];
  assign mem_29_2_W0_clk = W0_clk;
  assign mem_29_2_W0_data = W0_data[23:16];
  assign mem_29_2_W0_en = W0_en & W0_addr_sel == 8'h1d;
  assign mem_29_2_W0_mask = W0_mask[2];
  assign mem_29_3_R0_addr = R0_addr[25:0];
  assign mem_29_3_R0_clk = R0_clk;
  assign mem_29_3_R0_en = R0_en & R0_addr_sel == 8'h1d;
  assign mem_29_3_W0_addr = W0_addr[25:0];
  assign mem_29_3_W0_clk = W0_clk;
  assign mem_29_3_W0_data = W0_data[31:24];
  assign mem_29_3_W0_en = W0_en & W0_addr_sel == 8'h1d;
  assign mem_29_3_W0_mask = W0_mask[3];
  assign mem_29_4_R0_addr = R0_addr[25:0];
  assign mem_29_4_R0_clk = R0_clk;
  assign mem_29_4_R0_en = R0_en & R0_addr_sel == 8'h1d;
  assign mem_29_4_W0_addr = W0_addr[25:0];
  assign mem_29_4_W0_clk = W0_clk;
  assign mem_29_4_W0_data = W0_data[39:32];
  assign mem_29_4_W0_en = W0_en & W0_addr_sel == 8'h1d;
  assign mem_29_4_W0_mask = W0_mask[4];
  assign mem_29_5_R0_addr = R0_addr[25:0];
  assign mem_29_5_R0_clk = R0_clk;
  assign mem_29_5_R0_en = R0_en & R0_addr_sel == 8'h1d;
  assign mem_29_5_W0_addr = W0_addr[25:0];
  assign mem_29_5_W0_clk = W0_clk;
  assign mem_29_5_W0_data = W0_data[47:40];
  assign mem_29_5_W0_en = W0_en & W0_addr_sel == 8'h1d;
  assign mem_29_5_W0_mask = W0_mask[5];
  assign mem_29_6_R0_addr = R0_addr[25:0];
  assign mem_29_6_R0_clk = R0_clk;
  assign mem_29_6_R0_en = R0_en & R0_addr_sel == 8'h1d;
  assign mem_29_6_W0_addr = W0_addr[25:0];
  assign mem_29_6_W0_clk = W0_clk;
  assign mem_29_6_W0_data = W0_data[55:48];
  assign mem_29_6_W0_en = W0_en & W0_addr_sel == 8'h1d;
  assign mem_29_6_W0_mask = W0_mask[6];
  assign mem_29_7_R0_addr = R0_addr[25:0];
  assign mem_29_7_R0_clk = R0_clk;
  assign mem_29_7_R0_en = R0_en & R0_addr_sel == 8'h1d;
  assign mem_29_7_W0_addr = W0_addr[25:0];
  assign mem_29_7_W0_clk = W0_clk;
  assign mem_29_7_W0_data = W0_data[63:56];
  assign mem_29_7_W0_en = W0_en & W0_addr_sel == 8'h1d;
  assign mem_29_7_W0_mask = W0_mask[7];
  assign mem_30_0_R0_addr = R0_addr[25:0];
  assign mem_30_0_R0_clk = R0_clk;
  assign mem_30_0_R0_en = R0_en & R0_addr_sel == 8'h1e;
  assign mem_30_0_W0_addr = W0_addr[25:0];
  assign mem_30_0_W0_clk = W0_clk;
  assign mem_30_0_W0_data = W0_data[7:0];
  assign mem_30_0_W0_en = W0_en & W0_addr_sel == 8'h1e;
  assign mem_30_0_W0_mask = W0_mask[0];
  assign mem_30_1_R0_addr = R0_addr[25:0];
  assign mem_30_1_R0_clk = R0_clk;
  assign mem_30_1_R0_en = R0_en & R0_addr_sel == 8'h1e;
  assign mem_30_1_W0_addr = W0_addr[25:0];
  assign mem_30_1_W0_clk = W0_clk;
  assign mem_30_1_W0_data = W0_data[15:8];
  assign mem_30_1_W0_en = W0_en & W0_addr_sel == 8'h1e;
  assign mem_30_1_W0_mask = W0_mask[1];
  assign mem_30_2_R0_addr = R0_addr[25:0];
  assign mem_30_2_R0_clk = R0_clk;
  assign mem_30_2_R0_en = R0_en & R0_addr_sel == 8'h1e;
  assign mem_30_2_W0_addr = W0_addr[25:0];
  assign mem_30_2_W0_clk = W0_clk;
  assign mem_30_2_W0_data = W0_data[23:16];
  assign mem_30_2_W0_en = W0_en & W0_addr_sel == 8'h1e;
  assign mem_30_2_W0_mask = W0_mask[2];
  assign mem_30_3_R0_addr = R0_addr[25:0];
  assign mem_30_3_R0_clk = R0_clk;
  assign mem_30_3_R0_en = R0_en & R0_addr_sel == 8'h1e;
  assign mem_30_3_W0_addr = W0_addr[25:0];
  assign mem_30_3_W0_clk = W0_clk;
  assign mem_30_3_W0_data = W0_data[31:24];
  assign mem_30_3_W0_en = W0_en & W0_addr_sel == 8'h1e;
  assign mem_30_3_W0_mask = W0_mask[3];
  assign mem_30_4_R0_addr = R0_addr[25:0];
  assign mem_30_4_R0_clk = R0_clk;
  assign mem_30_4_R0_en = R0_en & R0_addr_sel == 8'h1e;
  assign mem_30_4_W0_addr = W0_addr[25:0];
  assign mem_30_4_W0_clk = W0_clk;
  assign mem_30_4_W0_data = W0_data[39:32];
  assign mem_30_4_W0_en = W0_en & W0_addr_sel == 8'h1e;
  assign mem_30_4_W0_mask = W0_mask[4];
  assign mem_30_5_R0_addr = R0_addr[25:0];
  assign mem_30_5_R0_clk = R0_clk;
  assign mem_30_5_R0_en = R0_en & R0_addr_sel == 8'h1e;
  assign mem_30_5_W0_addr = W0_addr[25:0];
  assign mem_30_5_W0_clk = W0_clk;
  assign mem_30_5_W0_data = W0_data[47:40];
  assign mem_30_5_W0_en = W0_en & W0_addr_sel == 8'h1e;
  assign mem_30_5_W0_mask = W0_mask[5];
  assign mem_30_6_R0_addr = R0_addr[25:0];
  assign mem_30_6_R0_clk = R0_clk;
  assign mem_30_6_R0_en = R0_en & R0_addr_sel == 8'h1e;
  assign mem_30_6_W0_addr = W0_addr[25:0];
  assign mem_30_6_W0_clk = W0_clk;
  assign mem_30_6_W0_data = W0_data[55:48];
  assign mem_30_6_W0_en = W0_en & W0_addr_sel == 8'h1e;
  assign mem_30_6_W0_mask = W0_mask[6];
  assign mem_30_7_R0_addr = R0_addr[25:0];
  assign mem_30_7_R0_clk = R0_clk;
  assign mem_30_7_R0_en = R0_en & R0_addr_sel == 8'h1e;
  assign mem_30_7_W0_addr = W0_addr[25:0];
  assign mem_30_7_W0_clk = W0_clk;
  assign mem_30_7_W0_data = W0_data[63:56];
  assign mem_30_7_W0_en = W0_en & W0_addr_sel == 8'h1e;
  assign mem_30_7_W0_mask = W0_mask[7];
  assign mem_31_0_R0_addr = R0_addr[25:0];
  assign mem_31_0_R0_clk = R0_clk;
  assign mem_31_0_R0_en = R0_en & R0_addr_sel == 8'h1f;
  assign mem_31_0_W0_addr = W0_addr[25:0];
  assign mem_31_0_W0_clk = W0_clk;
  assign mem_31_0_W0_data = W0_data[7:0];
  assign mem_31_0_W0_en = W0_en & W0_addr_sel == 8'h1f;
  assign mem_31_0_W0_mask = W0_mask[0];
  assign mem_31_1_R0_addr = R0_addr[25:0];
  assign mem_31_1_R0_clk = R0_clk;
  assign mem_31_1_R0_en = R0_en & R0_addr_sel == 8'h1f;
  assign mem_31_1_W0_addr = W0_addr[25:0];
  assign mem_31_1_W0_clk = W0_clk;
  assign mem_31_1_W0_data = W0_data[15:8];
  assign mem_31_1_W0_en = W0_en & W0_addr_sel == 8'h1f;
  assign mem_31_1_W0_mask = W0_mask[1];
  assign mem_31_2_R0_addr = R0_addr[25:0];
  assign mem_31_2_R0_clk = R0_clk;
  assign mem_31_2_R0_en = R0_en & R0_addr_sel == 8'h1f;
  assign mem_31_2_W0_addr = W0_addr[25:0];
  assign mem_31_2_W0_clk = W0_clk;
  assign mem_31_2_W0_data = W0_data[23:16];
  assign mem_31_2_W0_en = W0_en & W0_addr_sel == 8'h1f;
  assign mem_31_2_W0_mask = W0_mask[2];
  assign mem_31_3_R0_addr = R0_addr[25:0];
  assign mem_31_3_R0_clk = R0_clk;
  assign mem_31_3_R0_en = R0_en & R0_addr_sel == 8'h1f;
  assign mem_31_3_W0_addr = W0_addr[25:0];
  assign mem_31_3_W0_clk = W0_clk;
  assign mem_31_3_W0_data = W0_data[31:24];
  assign mem_31_3_W0_en = W0_en & W0_addr_sel == 8'h1f;
  assign mem_31_3_W0_mask = W0_mask[3];
  assign mem_31_4_R0_addr = R0_addr[25:0];
  assign mem_31_4_R0_clk = R0_clk;
  assign mem_31_4_R0_en = R0_en & R0_addr_sel == 8'h1f;
  assign mem_31_4_W0_addr = W0_addr[25:0];
  assign mem_31_4_W0_clk = W0_clk;
  assign mem_31_4_W0_data = W0_data[39:32];
  assign mem_31_4_W0_en = W0_en & W0_addr_sel == 8'h1f;
  assign mem_31_4_W0_mask = W0_mask[4];
  assign mem_31_5_R0_addr = R0_addr[25:0];
  assign mem_31_5_R0_clk = R0_clk;
  assign mem_31_5_R0_en = R0_en & R0_addr_sel == 8'h1f;
  assign mem_31_5_W0_addr = W0_addr[25:0];
  assign mem_31_5_W0_clk = W0_clk;
  assign mem_31_5_W0_data = W0_data[47:40];
  assign mem_31_5_W0_en = W0_en & W0_addr_sel == 8'h1f;
  assign mem_31_5_W0_mask = W0_mask[5];
  assign mem_31_6_R0_addr = R0_addr[25:0];
  assign mem_31_6_R0_clk = R0_clk;
  assign mem_31_6_R0_en = R0_en & R0_addr_sel == 8'h1f;
  assign mem_31_6_W0_addr = W0_addr[25:0];
  assign mem_31_6_W0_clk = W0_clk;
  assign mem_31_6_W0_data = W0_data[55:48];
  assign mem_31_6_W0_en = W0_en & W0_addr_sel == 8'h1f;
  assign mem_31_6_W0_mask = W0_mask[6];
  assign mem_31_7_R0_addr = R0_addr[25:0];
  assign mem_31_7_R0_clk = R0_clk;
  assign mem_31_7_R0_en = R0_en & R0_addr_sel == 8'h1f;
  assign mem_31_7_W0_addr = W0_addr[25:0];
  assign mem_31_7_W0_clk = W0_clk;
  assign mem_31_7_W0_data = W0_data[63:56];
  assign mem_31_7_W0_en = W0_en & W0_addr_sel == 8'h1f;
  assign mem_31_7_W0_mask = W0_mask[7];
  assign mem_32_0_R0_addr = R0_addr[25:0];
  assign mem_32_0_R0_clk = R0_clk;
  assign mem_32_0_R0_en = R0_en & R0_addr_sel == 8'h20;
  assign mem_32_0_W0_addr = W0_addr[25:0];
  assign mem_32_0_W0_clk = W0_clk;
  assign mem_32_0_W0_data = W0_data[7:0];
  assign mem_32_0_W0_en = W0_en & W0_addr_sel == 8'h20;
  assign mem_32_0_W0_mask = W0_mask[0];
  assign mem_32_1_R0_addr = R0_addr[25:0];
  assign mem_32_1_R0_clk = R0_clk;
  assign mem_32_1_R0_en = R0_en & R0_addr_sel == 8'h20;
  assign mem_32_1_W0_addr = W0_addr[25:0];
  assign mem_32_1_W0_clk = W0_clk;
  assign mem_32_1_W0_data = W0_data[15:8];
  assign mem_32_1_W0_en = W0_en & W0_addr_sel == 8'h20;
  assign mem_32_1_W0_mask = W0_mask[1];
  assign mem_32_2_R0_addr = R0_addr[25:0];
  assign mem_32_2_R0_clk = R0_clk;
  assign mem_32_2_R0_en = R0_en & R0_addr_sel == 8'h20;
  assign mem_32_2_W0_addr = W0_addr[25:0];
  assign mem_32_2_W0_clk = W0_clk;
  assign mem_32_2_W0_data = W0_data[23:16];
  assign mem_32_2_W0_en = W0_en & W0_addr_sel == 8'h20;
  assign mem_32_2_W0_mask = W0_mask[2];
  assign mem_32_3_R0_addr = R0_addr[25:0];
  assign mem_32_3_R0_clk = R0_clk;
  assign mem_32_3_R0_en = R0_en & R0_addr_sel == 8'h20;
  assign mem_32_3_W0_addr = W0_addr[25:0];
  assign mem_32_3_W0_clk = W0_clk;
  assign mem_32_3_W0_data = W0_data[31:24];
  assign mem_32_3_W0_en = W0_en & W0_addr_sel == 8'h20;
  assign mem_32_3_W0_mask = W0_mask[3];
  assign mem_32_4_R0_addr = R0_addr[25:0];
  assign mem_32_4_R0_clk = R0_clk;
  assign mem_32_4_R0_en = R0_en & R0_addr_sel == 8'h20;
  assign mem_32_4_W0_addr = W0_addr[25:0];
  assign mem_32_4_W0_clk = W0_clk;
  assign mem_32_4_W0_data = W0_data[39:32];
  assign mem_32_4_W0_en = W0_en & W0_addr_sel == 8'h20;
  assign mem_32_4_W0_mask = W0_mask[4];
  assign mem_32_5_R0_addr = R0_addr[25:0];
  assign mem_32_5_R0_clk = R0_clk;
  assign mem_32_5_R0_en = R0_en & R0_addr_sel == 8'h20;
  assign mem_32_5_W0_addr = W0_addr[25:0];
  assign mem_32_5_W0_clk = W0_clk;
  assign mem_32_5_W0_data = W0_data[47:40];
  assign mem_32_5_W0_en = W0_en & W0_addr_sel == 8'h20;
  assign mem_32_5_W0_mask = W0_mask[5];
  assign mem_32_6_R0_addr = R0_addr[25:0];
  assign mem_32_6_R0_clk = R0_clk;
  assign mem_32_6_R0_en = R0_en & R0_addr_sel == 8'h20;
  assign mem_32_6_W0_addr = W0_addr[25:0];
  assign mem_32_6_W0_clk = W0_clk;
  assign mem_32_6_W0_data = W0_data[55:48];
  assign mem_32_6_W0_en = W0_en & W0_addr_sel == 8'h20;
  assign mem_32_6_W0_mask = W0_mask[6];
  assign mem_32_7_R0_addr = R0_addr[25:0];
  assign mem_32_7_R0_clk = R0_clk;
  assign mem_32_7_R0_en = R0_en & R0_addr_sel == 8'h20;
  assign mem_32_7_W0_addr = W0_addr[25:0];
  assign mem_32_7_W0_clk = W0_clk;
  assign mem_32_7_W0_data = W0_data[63:56];
  assign mem_32_7_W0_en = W0_en & W0_addr_sel == 8'h20;
  assign mem_32_7_W0_mask = W0_mask[7];
  assign mem_33_0_R0_addr = R0_addr[25:0];
  assign mem_33_0_R0_clk = R0_clk;
  assign mem_33_0_R0_en = R0_en & R0_addr_sel == 8'h21;
  assign mem_33_0_W0_addr = W0_addr[25:0];
  assign mem_33_0_W0_clk = W0_clk;
  assign mem_33_0_W0_data = W0_data[7:0];
  assign mem_33_0_W0_en = W0_en & W0_addr_sel == 8'h21;
  assign mem_33_0_W0_mask = W0_mask[0];
  assign mem_33_1_R0_addr = R0_addr[25:0];
  assign mem_33_1_R0_clk = R0_clk;
  assign mem_33_1_R0_en = R0_en & R0_addr_sel == 8'h21;
  assign mem_33_1_W0_addr = W0_addr[25:0];
  assign mem_33_1_W0_clk = W0_clk;
  assign mem_33_1_W0_data = W0_data[15:8];
  assign mem_33_1_W0_en = W0_en & W0_addr_sel == 8'h21;
  assign mem_33_1_W0_mask = W0_mask[1];
  assign mem_33_2_R0_addr = R0_addr[25:0];
  assign mem_33_2_R0_clk = R0_clk;
  assign mem_33_2_R0_en = R0_en & R0_addr_sel == 8'h21;
  assign mem_33_2_W0_addr = W0_addr[25:0];
  assign mem_33_2_W0_clk = W0_clk;
  assign mem_33_2_W0_data = W0_data[23:16];
  assign mem_33_2_W0_en = W0_en & W0_addr_sel == 8'h21;
  assign mem_33_2_W0_mask = W0_mask[2];
  assign mem_33_3_R0_addr = R0_addr[25:0];
  assign mem_33_3_R0_clk = R0_clk;
  assign mem_33_3_R0_en = R0_en & R0_addr_sel == 8'h21;
  assign mem_33_3_W0_addr = W0_addr[25:0];
  assign mem_33_3_W0_clk = W0_clk;
  assign mem_33_3_W0_data = W0_data[31:24];
  assign mem_33_3_W0_en = W0_en & W0_addr_sel == 8'h21;
  assign mem_33_3_W0_mask = W0_mask[3];
  assign mem_33_4_R0_addr = R0_addr[25:0];
  assign mem_33_4_R0_clk = R0_clk;
  assign mem_33_4_R0_en = R0_en & R0_addr_sel == 8'h21;
  assign mem_33_4_W0_addr = W0_addr[25:0];
  assign mem_33_4_W0_clk = W0_clk;
  assign mem_33_4_W0_data = W0_data[39:32];
  assign mem_33_4_W0_en = W0_en & W0_addr_sel == 8'h21;
  assign mem_33_4_W0_mask = W0_mask[4];
  assign mem_33_5_R0_addr = R0_addr[25:0];
  assign mem_33_5_R0_clk = R0_clk;
  assign mem_33_5_R0_en = R0_en & R0_addr_sel == 8'h21;
  assign mem_33_5_W0_addr = W0_addr[25:0];
  assign mem_33_5_W0_clk = W0_clk;
  assign mem_33_5_W0_data = W0_data[47:40];
  assign mem_33_5_W0_en = W0_en & W0_addr_sel == 8'h21;
  assign mem_33_5_W0_mask = W0_mask[5];
  assign mem_33_6_R0_addr = R0_addr[25:0];
  assign mem_33_6_R0_clk = R0_clk;
  assign mem_33_6_R0_en = R0_en & R0_addr_sel == 8'h21;
  assign mem_33_6_W0_addr = W0_addr[25:0];
  assign mem_33_6_W0_clk = W0_clk;
  assign mem_33_6_W0_data = W0_data[55:48];
  assign mem_33_6_W0_en = W0_en & W0_addr_sel == 8'h21;
  assign mem_33_6_W0_mask = W0_mask[6];
  assign mem_33_7_R0_addr = R0_addr[25:0];
  assign mem_33_7_R0_clk = R0_clk;
  assign mem_33_7_R0_en = R0_en & R0_addr_sel == 8'h21;
  assign mem_33_7_W0_addr = W0_addr[25:0];
  assign mem_33_7_W0_clk = W0_clk;
  assign mem_33_7_W0_data = W0_data[63:56];
  assign mem_33_7_W0_en = W0_en & W0_addr_sel == 8'h21;
  assign mem_33_7_W0_mask = W0_mask[7];
  assign mem_34_0_R0_addr = R0_addr[25:0];
  assign mem_34_0_R0_clk = R0_clk;
  assign mem_34_0_R0_en = R0_en & R0_addr_sel == 8'h22;
  assign mem_34_0_W0_addr = W0_addr[25:0];
  assign mem_34_0_W0_clk = W0_clk;
  assign mem_34_0_W0_data = W0_data[7:0];
  assign mem_34_0_W0_en = W0_en & W0_addr_sel == 8'h22;
  assign mem_34_0_W0_mask = W0_mask[0];
  assign mem_34_1_R0_addr = R0_addr[25:0];
  assign mem_34_1_R0_clk = R0_clk;
  assign mem_34_1_R0_en = R0_en & R0_addr_sel == 8'h22;
  assign mem_34_1_W0_addr = W0_addr[25:0];
  assign mem_34_1_W0_clk = W0_clk;
  assign mem_34_1_W0_data = W0_data[15:8];
  assign mem_34_1_W0_en = W0_en & W0_addr_sel == 8'h22;
  assign mem_34_1_W0_mask = W0_mask[1];
  assign mem_34_2_R0_addr = R0_addr[25:0];
  assign mem_34_2_R0_clk = R0_clk;
  assign mem_34_2_R0_en = R0_en & R0_addr_sel == 8'h22;
  assign mem_34_2_W0_addr = W0_addr[25:0];
  assign mem_34_2_W0_clk = W0_clk;
  assign mem_34_2_W0_data = W0_data[23:16];
  assign mem_34_2_W0_en = W0_en & W0_addr_sel == 8'h22;
  assign mem_34_2_W0_mask = W0_mask[2];
  assign mem_34_3_R0_addr = R0_addr[25:0];
  assign mem_34_3_R0_clk = R0_clk;
  assign mem_34_3_R0_en = R0_en & R0_addr_sel == 8'h22;
  assign mem_34_3_W0_addr = W0_addr[25:0];
  assign mem_34_3_W0_clk = W0_clk;
  assign mem_34_3_W0_data = W0_data[31:24];
  assign mem_34_3_W0_en = W0_en & W0_addr_sel == 8'h22;
  assign mem_34_3_W0_mask = W0_mask[3];
  assign mem_34_4_R0_addr = R0_addr[25:0];
  assign mem_34_4_R0_clk = R0_clk;
  assign mem_34_4_R0_en = R0_en & R0_addr_sel == 8'h22;
  assign mem_34_4_W0_addr = W0_addr[25:0];
  assign mem_34_4_W0_clk = W0_clk;
  assign mem_34_4_W0_data = W0_data[39:32];
  assign mem_34_4_W0_en = W0_en & W0_addr_sel == 8'h22;
  assign mem_34_4_W0_mask = W0_mask[4];
  assign mem_34_5_R0_addr = R0_addr[25:0];
  assign mem_34_5_R0_clk = R0_clk;
  assign mem_34_5_R0_en = R0_en & R0_addr_sel == 8'h22;
  assign mem_34_5_W0_addr = W0_addr[25:0];
  assign mem_34_5_W0_clk = W0_clk;
  assign mem_34_5_W0_data = W0_data[47:40];
  assign mem_34_5_W0_en = W0_en & W0_addr_sel == 8'h22;
  assign mem_34_5_W0_mask = W0_mask[5];
  assign mem_34_6_R0_addr = R0_addr[25:0];
  assign mem_34_6_R0_clk = R0_clk;
  assign mem_34_6_R0_en = R0_en & R0_addr_sel == 8'h22;
  assign mem_34_6_W0_addr = W0_addr[25:0];
  assign mem_34_6_W0_clk = W0_clk;
  assign mem_34_6_W0_data = W0_data[55:48];
  assign mem_34_6_W0_en = W0_en & W0_addr_sel == 8'h22;
  assign mem_34_6_W0_mask = W0_mask[6];
  assign mem_34_7_R0_addr = R0_addr[25:0];
  assign mem_34_7_R0_clk = R0_clk;
  assign mem_34_7_R0_en = R0_en & R0_addr_sel == 8'h22;
  assign mem_34_7_W0_addr = W0_addr[25:0];
  assign mem_34_7_W0_clk = W0_clk;
  assign mem_34_7_W0_data = W0_data[63:56];
  assign mem_34_7_W0_en = W0_en & W0_addr_sel == 8'h22;
  assign mem_34_7_W0_mask = W0_mask[7];
  assign mem_35_0_R0_addr = R0_addr[25:0];
  assign mem_35_0_R0_clk = R0_clk;
  assign mem_35_0_R0_en = R0_en & R0_addr_sel == 8'h23;
  assign mem_35_0_W0_addr = W0_addr[25:0];
  assign mem_35_0_W0_clk = W0_clk;
  assign mem_35_0_W0_data = W0_data[7:0];
  assign mem_35_0_W0_en = W0_en & W0_addr_sel == 8'h23;
  assign mem_35_0_W0_mask = W0_mask[0];
  assign mem_35_1_R0_addr = R0_addr[25:0];
  assign mem_35_1_R0_clk = R0_clk;
  assign mem_35_1_R0_en = R0_en & R0_addr_sel == 8'h23;
  assign mem_35_1_W0_addr = W0_addr[25:0];
  assign mem_35_1_W0_clk = W0_clk;
  assign mem_35_1_W0_data = W0_data[15:8];
  assign mem_35_1_W0_en = W0_en & W0_addr_sel == 8'h23;
  assign mem_35_1_W0_mask = W0_mask[1];
  assign mem_35_2_R0_addr = R0_addr[25:0];
  assign mem_35_2_R0_clk = R0_clk;
  assign mem_35_2_R0_en = R0_en & R0_addr_sel == 8'h23;
  assign mem_35_2_W0_addr = W0_addr[25:0];
  assign mem_35_2_W0_clk = W0_clk;
  assign mem_35_2_W0_data = W0_data[23:16];
  assign mem_35_2_W0_en = W0_en & W0_addr_sel == 8'h23;
  assign mem_35_2_W0_mask = W0_mask[2];
  assign mem_35_3_R0_addr = R0_addr[25:0];
  assign mem_35_3_R0_clk = R0_clk;
  assign mem_35_3_R0_en = R0_en & R0_addr_sel == 8'h23;
  assign mem_35_3_W0_addr = W0_addr[25:0];
  assign mem_35_3_W0_clk = W0_clk;
  assign mem_35_3_W0_data = W0_data[31:24];
  assign mem_35_3_W0_en = W0_en & W0_addr_sel == 8'h23;
  assign mem_35_3_W0_mask = W0_mask[3];
  assign mem_35_4_R0_addr = R0_addr[25:0];
  assign mem_35_4_R0_clk = R0_clk;
  assign mem_35_4_R0_en = R0_en & R0_addr_sel == 8'h23;
  assign mem_35_4_W0_addr = W0_addr[25:0];
  assign mem_35_4_W0_clk = W0_clk;
  assign mem_35_4_W0_data = W0_data[39:32];
  assign mem_35_4_W0_en = W0_en & W0_addr_sel == 8'h23;
  assign mem_35_4_W0_mask = W0_mask[4];
  assign mem_35_5_R0_addr = R0_addr[25:0];
  assign mem_35_5_R0_clk = R0_clk;
  assign mem_35_5_R0_en = R0_en & R0_addr_sel == 8'h23;
  assign mem_35_5_W0_addr = W0_addr[25:0];
  assign mem_35_5_W0_clk = W0_clk;
  assign mem_35_5_W0_data = W0_data[47:40];
  assign mem_35_5_W0_en = W0_en & W0_addr_sel == 8'h23;
  assign mem_35_5_W0_mask = W0_mask[5];
  assign mem_35_6_R0_addr = R0_addr[25:0];
  assign mem_35_6_R0_clk = R0_clk;
  assign mem_35_6_R0_en = R0_en & R0_addr_sel == 8'h23;
  assign mem_35_6_W0_addr = W0_addr[25:0];
  assign mem_35_6_W0_clk = W0_clk;
  assign mem_35_6_W0_data = W0_data[55:48];
  assign mem_35_6_W0_en = W0_en & W0_addr_sel == 8'h23;
  assign mem_35_6_W0_mask = W0_mask[6];
  assign mem_35_7_R0_addr = R0_addr[25:0];
  assign mem_35_7_R0_clk = R0_clk;
  assign mem_35_7_R0_en = R0_en & R0_addr_sel == 8'h23;
  assign mem_35_7_W0_addr = W0_addr[25:0];
  assign mem_35_7_W0_clk = W0_clk;
  assign mem_35_7_W0_data = W0_data[63:56];
  assign mem_35_7_W0_en = W0_en & W0_addr_sel == 8'h23;
  assign mem_35_7_W0_mask = W0_mask[7];
  assign mem_36_0_R0_addr = R0_addr[25:0];
  assign mem_36_0_R0_clk = R0_clk;
  assign mem_36_0_R0_en = R0_en & R0_addr_sel == 8'h24;
  assign mem_36_0_W0_addr = W0_addr[25:0];
  assign mem_36_0_W0_clk = W0_clk;
  assign mem_36_0_W0_data = W0_data[7:0];
  assign mem_36_0_W0_en = W0_en & W0_addr_sel == 8'h24;
  assign mem_36_0_W0_mask = W0_mask[0];
  assign mem_36_1_R0_addr = R0_addr[25:0];
  assign mem_36_1_R0_clk = R0_clk;
  assign mem_36_1_R0_en = R0_en & R0_addr_sel == 8'h24;
  assign mem_36_1_W0_addr = W0_addr[25:0];
  assign mem_36_1_W0_clk = W0_clk;
  assign mem_36_1_W0_data = W0_data[15:8];
  assign mem_36_1_W0_en = W0_en & W0_addr_sel == 8'h24;
  assign mem_36_1_W0_mask = W0_mask[1];
  assign mem_36_2_R0_addr = R0_addr[25:0];
  assign mem_36_2_R0_clk = R0_clk;
  assign mem_36_2_R0_en = R0_en & R0_addr_sel == 8'h24;
  assign mem_36_2_W0_addr = W0_addr[25:0];
  assign mem_36_2_W0_clk = W0_clk;
  assign mem_36_2_W0_data = W0_data[23:16];
  assign mem_36_2_W0_en = W0_en & W0_addr_sel == 8'h24;
  assign mem_36_2_W0_mask = W0_mask[2];
  assign mem_36_3_R0_addr = R0_addr[25:0];
  assign mem_36_3_R0_clk = R0_clk;
  assign mem_36_3_R0_en = R0_en & R0_addr_sel == 8'h24;
  assign mem_36_3_W0_addr = W0_addr[25:0];
  assign mem_36_3_W0_clk = W0_clk;
  assign mem_36_3_W0_data = W0_data[31:24];
  assign mem_36_3_W0_en = W0_en & W0_addr_sel == 8'h24;
  assign mem_36_3_W0_mask = W0_mask[3];
  assign mem_36_4_R0_addr = R0_addr[25:0];
  assign mem_36_4_R0_clk = R0_clk;
  assign mem_36_4_R0_en = R0_en & R0_addr_sel == 8'h24;
  assign mem_36_4_W0_addr = W0_addr[25:0];
  assign mem_36_4_W0_clk = W0_clk;
  assign mem_36_4_W0_data = W0_data[39:32];
  assign mem_36_4_W0_en = W0_en & W0_addr_sel == 8'h24;
  assign mem_36_4_W0_mask = W0_mask[4];
  assign mem_36_5_R0_addr = R0_addr[25:0];
  assign mem_36_5_R0_clk = R0_clk;
  assign mem_36_5_R0_en = R0_en & R0_addr_sel == 8'h24;
  assign mem_36_5_W0_addr = W0_addr[25:0];
  assign mem_36_5_W0_clk = W0_clk;
  assign mem_36_5_W0_data = W0_data[47:40];
  assign mem_36_5_W0_en = W0_en & W0_addr_sel == 8'h24;
  assign mem_36_5_W0_mask = W0_mask[5];
  assign mem_36_6_R0_addr = R0_addr[25:0];
  assign mem_36_6_R0_clk = R0_clk;
  assign mem_36_6_R0_en = R0_en & R0_addr_sel == 8'h24;
  assign mem_36_6_W0_addr = W0_addr[25:0];
  assign mem_36_6_W0_clk = W0_clk;
  assign mem_36_6_W0_data = W0_data[55:48];
  assign mem_36_6_W0_en = W0_en & W0_addr_sel == 8'h24;
  assign mem_36_6_W0_mask = W0_mask[6];
  assign mem_36_7_R0_addr = R0_addr[25:0];
  assign mem_36_7_R0_clk = R0_clk;
  assign mem_36_7_R0_en = R0_en & R0_addr_sel == 8'h24;
  assign mem_36_7_W0_addr = W0_addr[25:0];
  assign mem_36_7_W0_clk = W0_clk;
  assign mem_36_7_W0_data = W0_data[63:56];
  assign mem_36_7_W0_en = W0_en & W0_addr_sel == 8'h24;
  assign mem_36_7_W0_mask = W0_mask[7];
  assign mem_37_0_R0_addr = R0_addr[25:0];
  assign mem_37_0_R0_clk = R0_clk;
  assign mem_37_0_R0_en = R0_en & R0_addr_sel == 8'h25;
  assign mem_37_0_W0_addr = W0_addr[25:0];
  assign mem_37_0_W0_clk = W0_clk;
  assign mem_37_0_W0_data = W0_data[7:0];
  assign mem_37_0_W0_en = W0_en & W0_addr_sel == 8'h25;
  assign mem_37_0_W0_mask = W0_mask[0];
  assign mem_37_1_R0_addr = R0_addr[25:0];
  assign mem_37_1_R0_clk = R0_clk;
  assign mem_37_1_R0_en = R0_en & R0_addr_sel == 8'h25;
  assign mem_37_1_W0_addr = W0_addr[25:0];
  assign mem_37_1_W0_clk = W0_clk;
  assign mem_37_1_W0_data = W0_data[15:8];
  assign mem_37_1_W0_en = W0_en & W0_addr_sel == 8'h25;
  assign mem_37_1_W0_mask = W0_mask[1];
  assign mem_37_2_R0_addr = R0_addr[25:0];
  assign mem_37_2_R0_clk = R0_clk;
  assign mem_37_2_R0_en = R0_en & R0_addr_sel == 8'h25;
  assign mem_37_2_W0_addr = W0_addr[25:0];
  assign mem_37_2_W0_clk = W0_clk;
  assign mem_37_2_W0_data = W0_data[23:16];
  assign mem_37_2_W0_en = W0_en & W0_addr_sel == 8'h25;
  assign mem_37_2_W0_mask = W0_mask[2];
  assign mem_37_3_R0_addr = R0_addr[25:0];
  assign mem_37_3_R0_clk = R0_clk;
  assign mem_37_3_R0_en = R0_en & R0_addr_sel == 8'h25;
  assign mem_37_3_W0_addr = W0_addr[25:0];
  assign mem_37_3_W0_clk = W0_clk;
  assign mem_37_3_W0_data = W0_data[31:24];
  assign mem_37_3_W0_en = W0_en & W0_addr_sel == 8'h25;
  assign mem_37_3_W0_mask = W0_mask[3];
  assign mem_37_4_R0_addr = R0_addr[25:0];
  assign mem_37_4_R0_clk = R0_clk;
  assign mem_37_4_R0_en = R0_en & R0_addr_sel == 8'h25;
  assign mem_37_4_W0_addr = W0_addr[25:0];
  assign mem_37_4_W0_clk = W0_clk;
  assign mem_37_4_W0_data = W0_data[39:32];
  assign mem_37_4_W0_en = W0_en & W0_addr_sel == 8'h25;
  assign mem_37_4_W0_mask = W0_mask[4];
  assign mem_37_5_R0_addr = R0_addr[25:0];
  assign mem_37_5_R0_clk = R0_clk;
  assign mem_37_5_R0_en = R0_en & R0_addr_sel == 8'h25;
  assign mem_37_5_W0_addr = W0_addr[25:0];
  assign mem_37_5_W0_clk = W0_clk;
  assign mem_37_5_W0_data = W0_data[47:40];
  assign mem_37_5_W0_en = W0_en & W0_addr_sel == 8'h25;
  assign mem_37_5_W0_mask = W0_mask[5];
  assign mem_37_6_R0_addr = R0_addr[25:0];
  assign mem_37_6_R0_clk = R0_clk;
  assign mem_37_6_R0_en = R0_en & R0_addr_sel == 8'h25;
  assign mem_37_6_W0_addr = W0_addr[25:0];
  assign mem_37_6_W0_clk = W0_clk;
  assign mem_37_6_W0_data = W0_data[55:48];
  assign mem_37_6_W0_en = W0_en & W0_addr_sel == 8'h25;
  assign mem_37_6_W0_mask = W0_mask[6];
  assign mem_37_7_R0_addr = R0_addr[25:0];
  assign mem_37_7_R0_clk = R0_clk;
  assign mem_37_7_R0_en = R0_en & R0_addr_sel == 8'h25;
  assign mem_37_7_W0_addr = W0_addr[25:0];
  assign mem_37_7_W0_clk = W0_clk;
  assign mem_37_7_W0_data = W0_data[63:56];
  assign mem_37_7_W0_en = W0_en & W0_addr_sel == 8'h25;
  assign mem_37_7_W0_mask = W0_mask[7];
  assign mem_38_0_R0_addr = R0_addr[25:0];
  assign mem_38_0_R0_clk = R0_clk;
  assign mem_38_0_R0_en = R0_en & R0_addr_sel == 8'h26;
  assign mem_38_0_W0_addr = W0_addr[25:0];
  assign mem_38_0_W0_clk = W0_clk;
  assign mem_38_0_W0_data = W0_data[7:0];
  assign mem_38_0_W0_en = W0_en & W0_addr_sel == 8'h26;
  assign mem_38_0_W0_mask = W0_mask[0];
  assign mem_38_1_R0_addr = R0_addr[25:0];
  assign mem_38_1_R0_clk = R0_clk;
  assign mem_38_1_R0_en = R0_en & R0_addr_sel == 8'h26;
  assign mem_38_1_W0_addr = W0_addr[25:0];
  assign mem_38_1_W0_clk = W0_clk;
  assign mem_38_1_W0_data = W0_data[15:8];
  assign mem_38_1_W0_en = W0_en & W0_addr_sel == 8'h26;
  assign mem_38_1_W0_mask = W0_mask[1];
  assign mem_38_2_R0_addr = R0_addr[25:0];
  assign mem_38_2_R0_clk = R0_clk;
  assign mem_38_2_R0_en = R0_en & R0_addr_sel == 8'h26;
  assign mem_38_2_W0_addr = W0_addr[25:0];
  assign mem_38_2_W0_clk = W0_clk;
  assign mem_38_2_W0_data = W0_data[23:16];
  assign mem_38_2_W0_en = W0_en & W0_addr_sel == 8'h26;
  assign mem_38_2_W0_mask = W0_mask[2];
  assign mem_38_3_R0_addr = R0_addr[25:0];
  assign mem_38_3_R0_clk = R0_clk;
  assign mem_38_3_R0_en = R0_en & R0_addr_sel == 8'h26;
  assign mem_38_3_W0_addr = W0_addr[25:0];
  assign mem_38_3_W0_clk = W0_clk;
  assign mem_38_3_W0_data = W0_data[31:24];
  assign mem_38_3_W0_en = W0_en & W0_addr_sel == 8'h26;
  assign mem_38_3_W0_mask = W0_mask[3];
  assign mem_38_4_R0_addr = R0_addr[25:0];
  assign mem_38_4_R0_clk = R0_clk;
  assign mem_38_4_R0_en = R0_en & R0_addr_sel == 8'h26;
  assign mem_38_4_W0_addr = W0_addr[25:0];
  assign mem_38_4_W0_clk = W0_clk;
  assign mem_38_4_W0_data = W0_data[39:32];
  assign mem_38_4_W0_en = W0_en & W0_addr_sel == 8'h26;
  assign mem_38_4_W0_mask = W0_mask[4];
  assign mem_38_5_R0_addr = R0_addr[25:0];
  assign mem_38_5_R0_clk = R0_clk;
  assign mem_38_5_R0_en = R0_en & R0_addr_sel == 8'h26;
  assign mem_38_5_W0_addr = W0_addr[25:0];
  assign mem_38_5_W0_clk = W0_clk;
  assign mem_38_5_W0_data = W0_data[47:40];
  assign mem_38_5_W0_en = W0_en & W0_addr_sel == 8'h26;
  assign mem_38_5_W0_mask = W0_mask[5];
  assign mem_38_6_R0_addr = R0_addr[25:0];
  assign mem_38_6_R0_clk = R0_clk;
  assign mem_38_6_R0_en = R0_en & R0_addr_sel == 8'h26;
  assign mem_38_6_W0_addr = W0_addr[25:0];
  assign mem_38_6_W0_clk = W0_clk;
  assign mem_38_6_W0_data = W0_data[55:48];
  assign mem_38_6_W0_en = W0_en & W0_addr_sel == 8'h26;
  assign mem_38_6_W0_mask = W0_mask[6];
  assign mem_38_7_R0_addr = R0_addr[25:0];
  assign mem_38_7_R0_clk = R0_clk;
  assign mem_38_7_R0_en = R0_en & R0_addr_sel == 8'h26;
  assign mem_38_7_W0_addr = W0_addr[25:0];
  assign mem_38_7_W0_clk = W0_clk;
  assign mem_38_7_W0_data = W0_data[63:56];
  assign mem_38_7_W0_en = W0_en & W0_addr_sel == 8'h26;
  assign mem_38_7_W0_mask = W0_mask[7];
  assign mem_39_0_R0_addr = R0_addr[25:0];
  assign mem_39_0_R0_clk = R0_clk;
  assign mem_39_0_R0_en = R0_en & R0_addr_sel == 8'h27;
  assign mem_39_0_W0_addr = W0_addr[25:0];
  assign mem_39_0_W0_clk = W0_clk;
  assign mem_39_0_W0_data = W0_data[7:0];
  assign mem_39_0_W0_en = W0_en & W0_addr_sel == 8'h27;
  assign mem_39_0_W0_mask = W0_mask[0];
  assign mem_39_1_R0_addr = R0_addr[25:0];
  assign mem_39_1_R0_clk = R0_clk;
  assign mem_39_1_R0_en = R0_en & R0_addr_sel == 8'h27;
  assign mem_39_1_W0_addr = W0_addr[25:0];
  assign mem_39_1_W0_clk = W0_clk;
  assign mem_39_1_W0_data = W0_data[15:8];
  assign mem_39_1_W0_en = W0_en & W0_addr_sel == 8'h27;
  assign mem_39_1_W0_mask = W0_mask[1];
  assign mem_39_2_R0_addr = R0_addr[25:0];
  assign mem_39_2_R0_clk = R0_clk;
  assign mem_39_2_R0_en = R0_en & R0_addr_sel == 8'h27;
  assign mem_39_2_W0_addr = W0_addr[25:0];
  assign mem_39_2_W0_clk = W0_clk;
  assign mem_39_2_W0_data = W0_data[23:16];
  assign mem_39_2_W0_en = W0_en & W0_addr_sel == 8'h27;
  assign mem_39_2_W0_mask = W0_mask[2];
  assign mem_39_3_R0_addr = R0_addr[25:0];
  assign mem_39_3_R0_clk = R0_clk;
  assign mem_39_3_R0_en = R0_en & R0_addr_sel == 8'h27;
  assign mem_39_3_W0_addr = W0_addr[25:0];
  assign mem_39_3_W0_clk = W0_clk;
  assign mem_39_3_W0_data = W0_data[31:24];
  assign mem_39_3_W0_en = W0_en & W0_addr_sel == 8'h27;
  assign mem_39_3_W0_mask = W0_mask[3];
  assign mem_39_4_R0_addr = R0_addr[25:0];
  assign mem_39_4_R0_clk = R0_clk;
  assign mem_39_4_R0_en = R0_en & R0_addr_sel == 8'h27;
  assign mem_39_4_W0_addr = W0_addr[25:0];
  assign mem_39_4_W0_clk = W0_clk;
  assign mem_39_4_W0_data = W0_data[39:32];
  assign mem_39_4_W0_en = W0_en & W0_addr_sel == 8'h27;
  assign mem_39_4_W0_mask = W0_mask[4];
  assign mem_39_5_R0_addr = R0_addr[25:0];
  assign mem_39_5_R0_clk = R0_clk;
  assign mem_39_5_R0_en = R0_en & R0_addr_sel == 8'h27;
  assign mem_39_5_W0_addr = W0_addr[25:0];
  assign mem_39_5_W0_clk = W0_clk;
  assign mem_39_5_W0_data = W0_data[47:40];
  assign mem_39_5_W0_en = W0_en & W0_addr_sel == 8'h27;
  assign mem_39_5_W0_mask = W0_mask[5];
  assign mem_39_6_R0_addr = R0_addr[25:0];
  assign mem_39_6_R0_clk = R0_clk;
  assign mem_39_6_R0_en = R0_en & R0_addr_sel == 8'h27;
  assign mem_39_6_W0_addr = W0_addr[25:0];
  assign mem_39_6_W0_clk = W0_clk;
  assign mem_39_6_W0_data = W0_data[55:48];
  assign mem_39_6_W0_en = W0_en & W0_addr_sel == 8'h27;
  assign mem_39_6_W0_mask = W0_mask[6];
  assign mem_39_7_R0_addr = R0_addr[25:0];
  assign mem_39_7_R0_clk = R0_clk;
  assign mem_39_7_R0_en = R0_en & R0_addr_sel == 8'h27;
  assign mem_39_7_W0_addr = W0_addr[25:0];
  assign mem_39_7_W0_clk = W0_clk;
  assign mem_39_7_W0_data = W0_data[63:56];
  assign mem_39_7_W0_en = W0_en & W0_addr_sel == 8'h27;
  assign mem_39_7_W0_mask = W0_mask[7];
  assign mem_40_0_R0_addr = R0_addr[25:0];
  assign mem_40_0_R0_clk = R0_clk;
  assign mem_40_0_R0_en = R0_en & R0_addr_sel == 8'h28;
  assign mem_40_0_W0_addr = W0_addr[25:0];
  assign mem_40_0_W0_clk = W0_clk;
  assign mem_40_0_W0_data = W0_data[7:0];
  assign mem_40_0_W0_en = W0_en & W0_addr_sel == 8'h28;
  assign mem_40_0_W0_mask = W0_mask[0];
  assign mem_40_1_R0_addr = R0_addr[25:0];
  assign mem_40_1_R0_clk = R0_clk;
  assign mem_40_1_R0_en = R0_en & R0_addr_sel == 8'h28;
  assign mem_40_1_W0_addr = W0_addr[25:0];
  assign mem_40_1_W0_clk = W0_clk;
  assign mem_40_1_W0_data = W0_data[15:8];
  assign mem_40_1_W0_en = W0_en & W0_addr_sel == 8'h28;
  assign mem_40_1_W0_mask = W0_mask[1];
  assign mem_40_2_R0_addr = R0_addr[25:0];
  assign mem_40_2_R0_clk = R0_clk;
  assign mem_40_2_R0_en = R0_en & R0_addr_sel == 8'h28;
  assign mem_40_2_W0_addr = W0_addr[25:0];
  assign mem_40_2_W0_clk = W0_clk;
  assign mem_40_2_W0_data = W0_data[23:16];
  assign mem_40_2_W0_en = W0_en & W0_addr_sel == 8'h28;
  assign mem_40_2_W0_mask = W0_mask[2];
  assign mem_40_3_R0_addr = R0_addr[25:0];
  assign mem_40_3_R0_clk = R0_clk;
  assign mem_40_3_R0_en = R0_en & R0_addr_sel == 8'h28;
  assign mem_40_3_W0_addr = W0_addr[25:0];
  assign mem_40_3_W0_clk = W0_clk;
  assign mem_40_3_W0_data = W0_data[31:24];
  assign mem_40_3_W0_en = W0_en & W0_addr_sel == 8'h28;
  assign mem_40_3_W0_mask = W0_mask[3];
  assign mem_40_4_R0_addr = R0_addr[25:0];
  assign mem_40_4_R0_clk = R0_clk;
  assign mem_40_4_R0_en = R0_en & R0_addr_sel == 8'h28;
  assign mem_40_4_W0_addr = W0_addr[25:0];
  assign mem_40_4_W0_clk = W0_clk;
  assign mem_40_4_W0_data = W0_data[39:32];
  assign mem_40_4_W0_en = W0_en & W0_addr_sel == 8'h28;
  assign mem_40_4_W0_mask = W0_mask[4];
  assign mem_40_5_R0_addr = R0_addr[25:0];
  assign mem_40_5_R0_clk = R0_clk;
  assign mem_40_5_R0_en = R0_en & R0_addr_sel == 8'h28;
  assign mem_40_5_W0_addr = W0_addr[25:0];
  assign mem_40_5_W0_clk = W0_clk;
  assign mem_40_5_W0_data = W0_data[47:40];
  assign mem_40_5_W0_en = W0_en & W0_addr_sel == 8'h28;
  assign mem_40_5_W0_mask = W0_mask[5];
  assign mem_40_6_R0_addr = R0_addr[25:0];
  assign mem_40_6_R0_clk = R0_clk;
  assign mem_40_6_R0_en = R0_en & R0_addr_sel == 8'h28;
  assign mem_40_6_W0_addr = W0_addr[25:0];
  assign mem_40_6_W0_clk = W0_clk;
  assign mem_40_6_W0_data = W0_data[55:48];
  assign mem_40_6_W0_en = W0_en & W0_addr_sel == 8'h28;
  assign mem_40_6_W0_mask = W0_mask[6];
  assign mem_40_7_R0_addr = R0_addr[25:0];
  assign mem_40_7_R0_clk = R0_clk;
  assign mem_40_7_R0_en = R0_en & R0_addr_sel == 8'h28;
  assign mem_40_7_W0_addr = W0_addr[25:0];
  assign mem_40_7_W0_clk = W0_clk;
  assign mem_40_7_W0_data = W0_data[63:56];
  assign mem_40_7_W0_en = W0_en & W0_addr_sel == 8'h28;
  assign mem_40_7_W0_mask = W0_mask[7];
  assign mem_41_0_R0_addr = R0_addr[25:0];
  assign mem_41_0_R0_clk = R0_clk;
  assign mem_41_0_R0_en = R0_en & R0_addr_sel == 8'h29;
  assign mem_41_0_W0_addr = W0_addr[25:0];
  assign mem_41_0_W0_clk = W0_clk;
  assign mem_41_0_W0_data = W0_data[7:0];
  assign mem_41_0_W0_en = W0_en & W0_addr_sel == 8'h29;
  assign mem_41_0_W0_mask = W0_mask[0];
  assign mem_41_1_R0_addr = R0_addr[25:0];
  assign mem_41_1_R0_clk = R0_clk;
  assign mem_41_1_R0_en = R0_en & R0_addr_sel == 8'h29;
  assign mem_41_1_W0_addr = W0_addr[25:0];
  assign mem_41_1_W0_clk = W0_clk;
  assign mem_41_1_W0_data = W0_data[15:8];
  assign mem_41_1_W0_en = W0_en & W0_addr_sel == 8'h29;
  assign mem_41_1_W0_mask = W0_mask[1];
  assign mem_41_2_R0_addr = R0_addr[25:0];
  assign mem_41_2_R0_clk = R0_clk;
  assign mem_41_2_R0_en = R0_en & R0_addr_sel == 8'h29;
  assign mem_41_2_W0_addr = W0_addr[25:0];
  assign mem_41_2_W0_clk = W0_clk;
  assign mem_41_2_W0_data = W0_data[23:16];
  assign mem_41_2_W0_en = W0_en & W0_addr_sel == 8'h29;
  assign mem_41_2_W0_mask = W0_mask[2];
  assign mem_41_3_R0_addr = R0_addr[25:0];
  assign mem_41_3_R0_clk = R0_clk;
  assign mem_41_3_R0_en = R0_en & R0_addr_sel == 8'h29;
  assign mem_41_3_W0_addr = W0_addr[25:0];
  assign mem_41_3_W0_clk = W0_clk;
  assign mem_41_3_W0_data = W0_data[31:24];
  assign mem_41_3_W0_en = W0_en & W0_addr_sel == 8'h29;
  assign mem_41_3_W0_mask = W0_mask[3];
  assign mem_41_4_R0_addr = R0_addr[25:0];
  assign mem_41_4_R0_clk = R0_clk;
  assign mem_41_4_R0_en = R0_en & R0_addr_sel == 8'h29;
  assign mem_41_4_W0_addr = W0_addr[25:0];
  assign mem_41_4_W0_clk = W0_clk;
  assign mem_41_4_W0_data = W0_data[39:32];
  assign mem_41_4_W0_en = W0_en & W0_addr_sel == 8'h29;
  assign mem_41_4_W0_mask = W0_mask[4];
  assign mem_41_5_R0_addr = R0_addr[25:0];
  assign mem_41_5_R0_clk = R0_clk;
  assign mem_41_5_R0_en = R0_en & R0_addr_sel == 8'h29;
  assign mem_41_5_W0_addr = W0_addr[25:0];
  assign mem_41_5_W0_clk = W0_clk;
  assign mem_41_5_W0_data = W0_data[47:40];
  assign mem_41_5_W0_en = W0_en & W0_addr_sel == 8'h29;
  assign mem_41_5_W0_mask = W0_mask[5];
  assign mem_41_6_R0_addr = R0_addr[25:0];
  assign mem_41_6_R0_clk = R0_clk;
  assign mem_41_6_R0_en = R0_en & R0_addr_sel == 8'h29;
  assign mem_41_6_W0_addr = W0_addr[25:0];
  assign mem_41_6_W0_clk = W0_clk;
  assign mem_41_6_W0_data = W0_data[55:48];
  assign mem_41_6_W0_en = W0_en & W0_addr_sel == 8'h29;
  assign mem_41_6_W0_mask = W0_mask[6];
  assign mem_41_7_R0_addr = R0_addr[25:0];
  assign mem_41_7_R0_clk = R0_clk;
  assign mem_41_7_R0_en = R0_en & R0_addr_sel == 8'h29;
  assign mem_41_7_W0_addr = W0_addr[25:0];
  assign mem_41_7_W0_clk = W0_clk;
  assign mem_41_7_W0_data = W0_data[63:56];
  assign mem_41_7_W0_en = W0_en & W0_addr_sel == 8'h29;
  assign mem_41_7_W0_mask = W0_mask[7];
  assign mem_42_0_R0_addr = R0_addr[25:0];
  assign mem_42_0_R0_clk = R0_clk;
  assign mem_42_0_R0_en = R0_en & R0_addr_sel == 8'h2a;
  assign mem_42_0_W0_addr = W0_addr[25:0];
  assign mem_42_0_W0_clk = W0_clk;
  assign mem_42_0_W0_data = W0_data[7:0];
  assign mem_42_0_W0_en = W0_en & W0_addr_sel == 8'h2a;
  assign mem_42_0_W0_mask = W0_mask[0];
  assign mem_42_1_R0_addr = R0_addr[25:0];
  assign mem_42_1_R0_clk = R0_clk;
  assign mem_42_1_R0_en = R0_en & R0_addr_sel == 8'h2a;
  assign mem_42_1_W0_addr = W0_addr[25:0];
  assign mem_42_1_W0_clk = W0_clk;
  assign mem_42_1_W0_data = W0_data[15:8];
  assign mem_42_1_W0_en = W0_en & W0_addr_sel == 8'h2a;
  assign mem_42_1_W0_mask = W0_mask[1];
  assign mem_42_2_R0_addr = R0_addr[25:0];
  assign mem_42_2_R0_clk = R0_clk;
  assign mem_42_2_R0_en = R0_en & R0_addr_sel == 8'h2a;
  assign mem_42_2_W0_addr = W0_addr[25:0];
  assign mem_42_2_W0_clk = W0_clk;
  assign mem_42_2_W0_data = W0_data[23:16];
  assign mem_42_2_W0_en = W0_en & W0_addr_sel == 8'h2a;
  assign mem_42_2_W0_mask = W0_mask[2];
  assign mem_42_3_R0_addr = R0_addr[25:0];
  assign mem_42_3_R0_clk = R0_clk;
  assign mem_42_3_R0_en = R0_en & R0_addr_sel == 8'h2a;
  assign mem_42_3_W0_addr = W0_addr[25:0];
  assign mem_42_3_W0_clk = W0_clk;
  assign mem_42_3_W0_data = W0_data[31:24];
  assign mem_42_3_W0_en = W0_en & W0_addr_sel == 8'h2a;
  assign mem_42_3_W0_mask = W0_mask[3];
  assign mem_42_4_R0_addr = R0_addr[25:0];
  assign mem_42_4_R0_clk = R0_clk;
  assign mem_42_4_R0_en = R0_en & R0_addr_sel == 8'h2a;
  assign mem_42_4_W0_addr = W0_addr[25:0];
  assign mem_42_4_W0_clk = W0_clk;
  assign mem_42_4_W0_data = W0_data[39:32];
  assign mem_42_4_W0_en = W0_en & W0_addr_sel == 8'h2a;
  assign mem_42_4_W0_mask = W0_mask[4];
  assign mem_42_5_R0_addr = R0_addr[25:0];
  assign mem_42_5_R0_clk = R0_clk;
  assign mem_42_5_R0_en = R0_en & R0_addr_sel == 8'h2a;
  assign mem_42_5_W0_addr = W0_addr[25:0];
  assign mem_42_5_W0_clk = W0_clk;
  assign mem_42_5_W0_data = W0_data[47:40];
  assign mem_42_5_W0_en = W0_en & W0_addr_sel == 8'h2a;
  assign mem_42_5_W0_mask = W0_mask[5];
  assign mem_42_6_R0_addr = R0_addr[25:0];
  assign mem_42_6_R0_clk = R0_clk;
  assign mem_42_6_R0_en = R0_en & R0_addr_sel == 8'h2a;
  assign mem_42_6_W0_addr = W0_addr[25:0];
  assign mem_42_6_W0_clk = W0_clk;
  assign mem_42_6_W0_data = W0_data[55:48];
  assign mem_42_6_W0_en = W0_en & W0_addr_sel == 8'h2a;
  assign mem_42_6_W0_mask = W0_mask[6];
  assign mem_42_7_R0_addr = R0_addr[25:0];
  assign mem_42_7_R0_clk = R0_clk;
  assign mem_42_7_R0_en = R0_en & R0_addr_sel == 8'h2a;
  assign mem_42_7_W0_addr = W0_addr[25:0];
  assign mem_42_7_W0_clk = W0_clk;
  assign mem_42_7_W0_data = W0_data[63:56];
  assign mem_42_7_W0_en = W0_en & W0_addr_sel == 8'h2a;
  assign mem_42_7_W0_mask = W0_mask[7];
  assign mem_43_0_R0_addr = R0_addr[25:0];
  assign mem_43_0_R0_clk = R0_clk;
  assign mem_43_0_R0_en = R0_en & R0_addr_sel == 8'h2b;
  assign mem_43_0_W0_addr = W0_addr[25:0];
  assign mem_43_0_W0_clk = W0_clk;
  assign mem_43_0_W0_data = W0_data[7:0];
  assign mem_43_0_W0_en = W0_en & W0_addr_sel == 8'h2b;
  assign mem_43_0_W0_mask = W0_mask[0];
  assign mem_43_1_R0_addr = R0_addr[25:0];
  assign mem_43_1_R0_clk = R0_clk;
  assign mem_43_1_R0_en = R0_en & R0_addr_sel == 8'h2b;
  assign mem_43_1_W0_addr = W0_addr[25:0];
  assign mem_43_1_W0_clk = W0_clk;
  assign mem_43_1_W0_data = W0_data[15:8];
  assign mem_43_1_W0_en = W0_en & W0_addr_sel == 8'h2b;
  assign mem_43_1_W0_mask = W0_mask[1];
  assign mem_43_2_R0_addr = R0_addr[25:0];
  assign mem_43_2_R0_clk = R0_clk;
  assign mem_43_2_R0_en = R0_en & R0_addr_sel == 8'h2b;
  assign mem_43_2_W0_addr = W0_addr[25:0];
  assign mem_43_2_W0_clk = W0_clk;
  assign mem_43_2_W0_data = W0_data[23:16];
  assign mem_43_2_W0_en = W0_en & W0_addr_sel == 8'h2b;
  assign mem_43_2_W0_mask = W0_mask[2];
  assign mem_43_3_R0_addr = R0_addr[25:0];
  assign mem_43_3_R0_clk = R0_clk;
  assign mem_43_3_R0_en = R0_en & R0_addr_sel == 8'h2b;
  assign mem_43_3_W0_addr = W0_addr[25:0];
  assign mem_43_3_W0_clk = W0_clk;
  assign mem_43_3_W0_data = W0_data[31:24];
  assign mem_43_3_W0_en = W0_en & W0_addr_sel == 8'h2b;
  assign mem_43_3_W0_mask = W0_mask[3];
  assign mem_43_4_R0_addr = R0_addr[25:0];
  assign mem_43_4_R0_clk = R0_clk;
  assign mem_43_4_R0_en = R0_en & R0_addr_sel == 8'h2b;
  assign mem_43_4_W0_addr = W0_addr[25:0];
  assign mem_43_4_W0_clk = W0_clk;
  assign mem_43_4_W0_data = W0_data[39:32];
  assign mem_43_4_W0_en = W0_en & W0_addr_sel == 8'h2b;
  assign mem_43_4_W0_mask = W0_mask[4];
  assign mem_43_5_R0_addr = R0_addr[25:0];
  assign mem_43_5_R0_clk = R0_clk;
  assign mem_43_5_R0_en = R0_en & R0_addr_sel == 8'h2b;
  assign mem_43_5_W0_addr = W0_addr[25:0];
  assign mem_43_5_W0_clk = W0_clk;
  assign mem_43_5_W0_data = W0_data[47:40];
  assign mem_43_5_W0_en = W0_en & W0_addr_sel == 8'h2b;
  assign mem_43_5_W0_mask = W0_mask[5];
  assign mem_43_6_R0_addr = R0_addr[25:0];
  assign mem_43_6_R0_clk = R0_clk;
  assign mem_43_6_R0_en = R0_en & R0_addr_sel == 8'h2b;
  assign mem_43_6_W0_addr = W0_addr[25:0];
  assign mem_43_6_W0_clk = W0_clk;
  assign mem_43_6_W0_data = W0_data[55:48];
  assign mem_43_6_W0_en = W0_en & W0_addr_sel == 8'h2b;
  assign mem_43_6_W0_mask = W0_mask[6];
  assign mem_43_7_R0_addr = R0_addr[25:0];
  assign mem_43_7_R0_clk = R0_clk;
  assign mem_43_7_R0_en = R0_en & R0_addr_sel == 8'h2b;
  assign mem_43_7_W0_addr = W0_addr[25:0];
  assign mem_43_7_W0_clk = W0_clk;
  assign mem_43_7_W0_data = W0_data[63:56];
  assign mem_43_7_W0_en = W0_en & W0_addr_sel == 8'h2b;
  assign mem_43_7_W0_mask = W0_mask[7];
  assign mem_44_0_R0_addr = R0_addr[25:0];
  assign mem_44_0_R0_clk = R0_clk;
  assign mem_44_0_R0_en = R0_en & R0_addr_sel == 8'h2c;
  assign mem_44_0_W0_addr = W0_addr[25:0];
  assign mem_44_0_W0_clk = W0_clk;
  assign mem_44_0_W0_data = W0_data[7:0];
  assign mem_44_0_W0_en = W0_en & W0_addr_sel == 8'h2c;
  assign mem_44_0_W0_mask = W0_mask[0];
  assign mem_44_1_R0_addr = R0_addr[25:0];
  assign mem_44_1_R0_clk = R0_clk;
  assign mem_44_1_R0_en = R0_en & R0_addr_sel == 8'h2c;
  assign mem_44_1_W0_addr = W0_addr[25:0];
  assign mem_44_1_W0_clk = W0_clk;
  assign mem_44_1_W0_data = W0_data[15:8];
  assign mem_44_1_W0_en = W0_en & W0_addr_sel == 8'h2c;
  assign mem_44_1_W0_mask = W0_mask[1];
  assign mem_44_2_R0_addr = R0_addr[25:0];
  assign mem_44_2_R0_clk = R0_clk;
  assign mem_44_2_R0_en = R0_en & R0_addr_sel == 8'h2c;
  assign mem_44_2_W0_addr = W0_addr[25:0];
  assign mem_44_2_W0_clk = W0_clk;
  assign mem_44_2_W0_data = W0_data[23:16];
  assign mem_44_2_W0_en = W0_en & W0_addr_sel == 8'h2c;
  assign mem_44_2_W0_mask = W0_mask[2];
  assign mem_44_3_R0_addr = R0_addr[25:0];
  assign mem_44_3_R0_clk = R0_clk;
  assign mem_44_3_R0_en = R0_en & R0_addr_sel == 8'h2c;
  assign mem_44_3_W0_addr = W0_addr[25:0];
  assign mem_44_3_W0_clk = W0_clk;
  assign mem_44_3_W0_data = W0_data[31:24];
  assign mem_44_3_W0_en = W0_en & W0_addr_sel == 8'h2c;
  assign mem_44_3_W0_mask = W0_mask[3];
  assign mem_44_4_R0_addr = R0_addr[25:0];
  assign mem_44_4_R0_clk = R0_clk;
  assign mem_44_4_R0_en = R0_en & R0_addr_sel == 8'h2c;
  assign mem_44_4_W0_addr = W0_addr[25:0];
  assign mem_44_4_W0_clk = W0_clk;
  assign mem_44_4_W0_data = W0_data[39:32];
  assign mem_44_4_W0_en = W0_en & W0_addr_sel == 8'h2c;
  assign mem_44_4_W0_mask = W0_mask[4];
  assign mem_44_5_R0_addr = R0_addr[25:0];
  assign mem_44_5_R0_clk = R0_clk;
  assign mem_44_5_R0_en = R0_en & R0_addr_sel == 8'h2c;
  assign mem_44_5_W0_addr = W0_addr[25:0];
  assign mem_44_5_W0_clk = W0_clk;
  assign mem_44_5_W0_data = W0_data[47:40];
  assign mem_44_5_W0_en = W0_en & W0_addr_sel == 8'h2c;
  assign mem_44_5_W0_mask = W0_mask[5];
  assign mem_44_6_R0_addr = R0_addr[25:0];
  assign mem_44_6_R0_clk = R0_clk;
  assign mem_44_6_R0_en = R0_en & R0_addr_sel == 8'h2c;
  assign mem_44_6_W0_addr = W0_addr[25:0];
  assign mem_44_6_W0_clk = W0_clk;
  assign mem_44_6_W0_data = W0_data[55:48];
  assign mem_44_6_W0_en = W0_en & W0_addr_sel == 8'h2c;
  assign mem_44_6_W0_mask = W0_mask[6];
  assign mem_44_7_R0_addr = R0_addr[25:0];
  assign mem_44_7_R0_clk = R0_clk;
  assign mem_44_7_R0_en = R0_en & R0_addr_sel == 8'h2c;
  assign mem_44_7_W0_addr = W0_addr[25:0];
  assign mem_44_7_W0_clk = W0_clk;
  assign mem_44_7_W0_data = W0_data[63:56];
  assign mem_44_7_W0_en = W0_en & W0_addr_sel == 8'h2c;
  assign mem_44_7_W0_mask = W0_mask[7];
  assign mem_45_0_R0_addr = R0_addr[25:0];
  assign mem_45_0_R0_clk = R0_clk;
  assign mem_45_0_R0_en = R0_en & R0_addr_sel == 8'h2d;
  assign mem_45_0_W0_addr = W0_addr[25:0];
  assign mem_45_0_W0_clk = W0_clk;
  assign mem_45_0_W0_data = W0_data[7:0];
  assign mem_45_0_W0_en = W0_en & W0_addr_sel == 8'h2d;
  assign mem_45_0_W0_mask = W0_mask[0];
  assign mem_45_1_R0_addr = R0_addr[25:0];
  assign mem_45_1_R0_clk = R0_clk;
  assign mem_45_1_R0_en = R0_en & R0_addr_sel == 8'h2d;
  assign mem_45_1_W0_addr = W0_addr[25:0];
  assign mem_45_1_W0_clk = W0_clk;
  assign mem_45_1_W0_data = W0_data[15:8];
  assign mem_45_1_W0_en = W0_en & W0_addr_sel == 8'h2d;
  assign mem_45_1_W0_mask = W0_mask[1];
  assign mem_45_2_R0_addr = R0_addr[25:0];
  assign mem_45_2_R0_clk = R0_clk;
  assign mem_45_2_R0_en = R0_en & R0_addr_sel == 8'h2d;
  assign mem_45_2_W0_addr = W0_addr[25:0];
  assign mem_45_2_W0_clk = W0_clk;
  assign mem_45_2_W0_data = W0_data[23:16];
  assign mem_45_2_W0_en = W0_en & W0_addr_sel == 8'h2d;
  assign mem_45_2_W0_mask = W0_mask[2];
  assign mem_45_3_R0_addr = R0_addr[25:0];
  assign mem_45_3_R0_clk = R0_clk;
  assign mem_45_3_R0_en = R0_en & R0_addr_sel == 8'h2d;
  assign mem_45_3_W0_addr = W0_addr[25:0];
  assign mem_45_3_W0_clk = W0_clk;
  assign mem_45_3_W0_data = W0_data[31:24];
  assign mem_45_3_W0_en = W0_en & W0_addr_sel == 8'h2d;
  assign mem_45_3_W0_mask = W0_mask[3];
  assign mem_45_4_R0_addr = R0_addr[25:0];
  assign mem_45_4_R0_clk = R0_clk;
  assign mem_45_4_R0_en = R0_en & R0_addr_sel == 8'h2d;
  assign mem_45_4_W0_addr = W0_addr[25:0];
  assign mem_45_4_W0_clk = W0_clk;
  assign mem_45_4_W0_data = W0_data[39:32];
  assign mem_45_4_W0_en = W0_en & W0_addr_sel == 8'h2d;
  assign mem_45_4_W0_mask = W0_mask[4];
  assign mem_45_5_R0_addr = R0_addr[25:0];
  assign mem_45_5_R0_clk = R0_clk;
  assign mem_45_5_R0_en = R0_en & R0_addr_sel == 8'h2d;
  assign mem_45_5_W0_addr = W0_addr[25:0];
  assign mem_45_5_W0_clk = W0_clk;
  assign mem_45_5_W0_data = W0_data[47:40];
  assign mem_45_5_W0_en = W0_en & W0_addr_sel == 8'h2d;
  assign mem_45_5_W0_mask = W0_mask[5];
  assign mem_45_6_R0_addr = R0_addr[25:0];
  assign mem_45_6_R0_clk = R0_clk;
  assign mem_45_6_R0_en = R0_en & R0_addr_sel == 8'h2d;
  assign mem_45_6_W0_addr = W0_addr[25:0];
  assign mem_45_6_W0_clk = W0_clk;
  assign mem_45_6_W0_data = W0_data[55:48];
  assign mem_45_6_W0_en = W0_en & W0_addr_sel == 8'h2d;
  assign mem_45_6_W0_mask = W0_mask[6];
  assign mem_45_7_R0_addr = R0_addr[25:0];
  assign mem_45_7_R0_clk = R0_clk;
  assign mem_45_7_R0_en = R0_en & R0_addr_sel == 8'h2d;
  assign mem_45_7_W0_addr = W0_addr[25:0];
  assign mem_45_7_W0_clk = W0_clk;
  assign mem_45_7_W0_data = W0_data[63:56];
  assign mem_45_7_W0_en = W0_en & W0_addr_sel == 8'h2d;
  assign mem_45_7_W0_mask = W0_mask[7];
  assign mem_46_0_R0_addr = R0_addr[25:0];
  assign mem_46_0_R0_clk = R0_clk;
  assign mem_46_0_R0_en = R0_en & R0_addr_sel == 8'h2e;
  assign mem_46_0_W0_addr = W0_addr[25:0];
  assign mem_46_0_W0_clk = W0_clk;
  assign mem_46_0_W0_data = W0_data[7:0];
  assign mem_46_0_W0_en = W0_en & W0_addr_sel == 8'h2e;
  assign mem_46_0_W0_mask = W0_mask[0];
  assign mem_46_1_R0_addr = R0_addr[25:0];
  assign mem_46_1_R0_clk = R0_clk;
  assign mem_46_1_R0_en = R0_en & R0_addr_sel == 8'h2e;
  assign mem_46_1_W0_addr = W0_addr[25:0];
  assign mem_46_1_W0_clk = W0_clk;
  assign mem_46_1_W0_data = W0_data[15:8];
  assign mem_46_1_W0_en = W0_en & W0_addr_sel == 8'h2e;
  assign mem_46_1_W0_mask = W0_mask[1];
  assign mem_46_2_R0_addr = R0_addr[25:0];
  assign mem_46_2_R0_clk = R0_clk;
  assign mem_46_2_R0_en = R0_en & R0_addr_sel == 8'h2e;
  assign mem_46_2_W0_addr = W0_addr[25:0];
  assign mem_46_2_W0_clk = W0_clk;
  assign mem_46_2_W0_data = W0_data[23:16];
  assign mem_46_2_W0_en = W0_en & W0_addr_sel == 8'h2e;
  assign mem_46_2_W0_mask = W0_mask[2];
  assign mem_46_3_R0_addr = R0_addr[25:0];
  assign mem_46_3_R0_clk = R0_clk;
  assign mem_46_3_R0_en = R0_en & R0_addr_sel == 8'h2e;
  assign mem_46_3_W0_addr = W0_addr[25:0];
  assign mem_46_3_W0_clk = W0_clk;
  assign mem_46_3_W0_data = W0_data[31:24];
  assign mem_46_3_W0_en = W0_en & W0_addr_sel == 8'h2e;
  assign mem_46_3_W0_mask = W0_mask[3];
  assign mem_46_4_R0_addr = R0_addr[25:0];
  assign mem_46_4_R0_clk = R0_clk;
  assign mem_46_4_R0_en = R0_en & R0_addr_sel == 8'h2e;
  assign mem_46_4_W0_addr = W0_addr[25:0];
  assign mem_46_4_W0_clk = W0_clk;
  assign mem_46_4_W0_data = W0_data[39:32];
  assign mem_46_4_W0_en = W0_en & W0_addr_sel == 8'h2e;
  assign mem_46_4_W0_mask = W0_mask[4];
  assign mem_46_5_R0_addr = R0_addr[25:0];
  assign mem_46_5_R0_clk = R0_clk;
  assign mem_46_5_R0_en = R0_en & R0_addr_sel == 8'h2e;
  assign mem_46_5_W0_addr = W0_addr[25:0];
  assign mem_46_5_W0_clk = W0_clk;
  assign mem_46_5_W0_data = W0_data[47:40];
  assign mem_46_5_W0_en = W0_en & W0_addr_sel == 8'h2e;
  assign mem_46_5_W0_mask = W0_mask[5];
  assign mem_46_6_R0_addr = R0_addr[25:0];
  assign mem_46_6_R0_clk = R0_clk;
  assign mem_46_6_R0_en = R0_en & R0_addr_sel == 8'h2e;
  assign mem_46_6_W0_addr = W0_addr[25:0];
  assign mem_46_6_W0_clk = W0_clk;
  assign mem_46_6_W0_data = W0_data[55:48];
  assign mem_46_6_W0_en = W0_en & W0_addr_sel == 8'h2e;
  assign mem_46_6_W0_mask = W0_mask[6];
  assign mem_46_7_R0_addr = R0_addr[25:0];
  assign mem_46_7_R0_clk = R0_clk;
  assign mem_46_7_R0_en = R0_en & R0_addr_sel == 8'h2e;
  assign mem_46_7_W0_addr = W0_addr[25:0];
  assign mem_46_7_W0_clk = W0_clk;
  assign mem_46_7_W0_data = W0_data[63:56];
  assign mem_46_7_W0_en = W0_en & W0_addr_sel == 8'h2e;
  assign mem_46_7_W0_mask = W0_mask[7];
  assign mem_47_0_R0_addr = R0_addr[25:0];
  assign mem_47_0_R0_clk = R0_clk;
  assign mem_47_0_R0_en = R0_en & R0_addr_sel == 8'h2f;
  assign mem_47_0_W0_addr = W0_addr[25:0];
  assign mem_47_0_W0_clk = W0_clk;
  assign mem_47_0_W0_data = W0_data[7:0];
  assign mem_47_0_W0_en = W0_en & W0_addr_sel == 8'h2f;
  assign mem_47_0_W0_mask = W0_mask[0];
  assign mem_47_1_R0_addr = R0_addr[25:0];
  assign mem_47_1_R0_clk = R0_clk;
  assign mem_47_1_R0_en = R0_en & R0_addr_sel == 8'h2f;
  assign mem_47_1_W0_addr = W0_addr[25:0];
  assign mem_47_1_W0_clk = W0_clk;
  assign mem_47_1_W0_data = W0_data[15:8];
  assign mem_47_1_W0_en = W0_en & W0_addr_sel == 8'h2f;
  assign mem_47_1_W0_mask = W0_mask[1];
  assign mem_47_2_R0_addr = R0_addr[25:0];
  assign mem_47_2_R0_clk = R0_clk;
  assign mem_47_2_R0_en = R0_en & R0_addr_sel == 8'h2f;
  assign mem_47_2_W0_addr = W0_addr[25:0];
  assign mem_47_2_W0_clk = W0_clk;
  assign mem_47_2_W0_data = W0_data[23:16];
  assign mem_47_2_W0_en = W0_en & W0_addr_sel == 8'h2f;
  assign mem_47_2_W0_mask = W0_mask[2];
  assign mem_47_3_R0_addr = R0_addr[25:0];
  assign mem_47_3_R0_clk = R0_clk;
  assign mem_47_3_R0_en = R0_en & R0_addr_sel == 8'h2f;
  assign mem_47_3_W0_addr = W0_addr[25:0];
  assign mem_47_3_W0_clk = W0_clk;
  assign mem_47_3_W0_data = W0_data[31:24];
  assign mem_47_3_W0_en = W0_en & W0_addr_sel == 8'h2f;
  assign mem_47_3_W0_mask = W0_mask[3];
  assign mem_47_4_R0_addr = R0_addr[25:0];
  assign mem_47_4_R0_clk = R0_clk;
  assign mem_47_4_R0_en = R0_en & R0_addr_sel == 8'h2f;
  assign mem_47_4_W0_addr = W0_addr[25:0];
  assign mem_47_4_W0_clk = W0_clk;
  assign mem_47_4_W0_data = W0_data[39:32];
  assign mem_47_4_W0_en = W0_en & W0_addr_sel == 8'h2f;
  assign mem_47_4_W0_mask = W0_mask[4];
  assign mem_47_5_R0_addr = R0_addr[25:0];
  assign mem_47_5_R0_clk = R0_clk;
  assign mem_47_5_R0_en = R0_en & R0_addr_sel == 8'h2f;
  assign mem_47_5_W0_addr = W0_addr[25:0];
  assign mem_47_5_W0_clk = W0_clk;
  assign mem_47_5_W0_data = W0_data[47:40];
  assign mem_47_5_W0_en = W0_en & W0_addr_sel == 8'h2f;
  assign mem_47_5_W0_mask = W0_mask[5];
  assign mem_47_6_R0_addr = R0_addr[25:0];
  assign mem_47_6_R0_clk = R0_clk;
  assign mem_47_6_R0_en = R0_en & R0_addr_sel == 8'h2f;
  assign mem_47_6_W0_addr = W0_addr[25:0];
  assign mem_47_6_W0_clk = W0_clk;
  assign mem_47_6_W0_data = W0_data[55:48];
  assign mem_47_6_W0_en = W0_en & W0_addr_sel == 8'h2f;
  assign mem_47_6_W0_mask = W0_mask[6];
  assign mem_47_7_R0_addr = R0_addr[25:0];
  assign mem_47_7_R0_clk = R0_clk;
  assign mem_47_7_R0_en = R0_en & R0_addr_sel == 8'h2f;
  assign mem_47_7_W0_addr = W0_addr[25:0];
  assign mem_47_7_W0_clk = W0_clk;
  assign mem_47_7_W0_data = W0_data[63:56];
  assign mem_47_7_W0_en = W0_en & W0_addr_sel == 8'h2f;
  assign mem_47_7_W0_mask = W0_mask[7];
  assign mem_48_0_R0_addr = R0_addr[25:0];
  assign mem_48_0_R0_clk = R0_clk;
  assign mem_48_0_R0_en = R0_en & R0_addr_sel == 8'h30;
  assign mem_48_0_W0_addr = W0_addr[25:0];
  assign mem_48_0_W0_clk = W0_clk;
  assign mem_48_0_W0_data = W0_data[7:0];
  assign mem_48_0_W0_en = W0_en & W0_addr_sel == 8'h30;
  assign mem_48_0_W0_mask = W0_mask[0];
  assign mem_48_1_R0_addr = R0_addr[25:0];
  assign mem_48_1_R0_clk = R0_clk;
  assign mem_48_1_R0_en = R0_en & R0_addr_sel == 8'h30;
  assign mem_48_1_W0_addr = W0_addr[25:0];
  assign mem_48_1_W0_clk = W0_clk;
  assign mem_48_1_W0_data = W0_data[15:8];
  assign mem_48_1_W0_en = W0_en & W0_addr_sel == 8'h30;
  assign mem_48_1_W0_mask = W0_mask[1];
  assign mem_48_2_R0_addr = R0_addr[25:0];
  assign mem_48_2_R0_clk = R0_clk;
  assign mem_48_2_R0_en = R0_en & R0_addr_sel == 8'h30;
  assign mem_48_2_W0_addr = W0_addr[25:0];
  assign mem_48_2_W0_clk = W0_clk;
  assign mem_48_2_W0_data = W0_data[23:16];
  assign mem_48_2_W0_en = W0_en & W0_addr_sel == 8'h30;
  assign mem_48_2_W0_mask = W0_mask[2];
  assign mem_48_3_R0_addr = R0_addr[25:0];
  assign mem_48_3_R0_clk = R0_clk;
  assign mem_48_3_R0_en = R0_en & R0_addr_sel == 8'h30;
  assign mem_48_3_W0_addr = W0_addr[25:0];
  assign mem_48_3_W0_clk = W0_clk;
  assign mem_48_3_W0_data = W0_data[31:24];
  assign mem_48_3_W0_en = W0_en & W0_addr_sel == 8'h30;
  assign mem_48_3_W0_mask = W0_mask[3];
  assign mem_48_4_R0_addr = R0_addr[25:0];
  assign mem_48_4_R0_clk = R0_clk;
  assign mem_48_4_R0_en = R0_en & R0_addr_sel == 8'h30;
  assign mem_48_4_W0_addr = W0_addr[25:0];
  assign mem_48_4_W0_clk = W0_clk;
  assign mem_48_4_W0_data = W0_data[39:32];
  assign mem_48_4_W0_en = W0_en & W0_addr_sel == 8'h30;
  assign mem_48_4_W0_mask = W0_mask[4];
  assign mem_48_5_R0_addr = R0_addr[25:0];
  assign mem_48_5_R0_clk = R0_clk;
  assign mem_48_5_R0_en = R0_en & R0_addr_sel == 8'h30;
  assign mem_48_5_W0_addr = W0_addr[25:0];
  assign mem_48_5_W0_clk = W0_clk;
  assign mem_48_5_W0_data = W0_data[47:40];
  assign mem_48_5_W0_en = W0_en & W0_addr_sel == 8'h30;
  assign mem_48_5_W0_mask = W0_mask[5];
  assign mem_48_6_R0_addr = R0_addr[25:0];
  assign mem_48_6_R0_clk = R0_clk;
  assign mem_48_6_R0_en = R0_en & R0_addr_sel == 8'h30;
  assign mem_48_6_W0_addr = W0_addr[25:0];
  assign mem_48_6_W0_clk = W0_clk;
  assign mem_48_6_W0_data = W0_data[55:48];
  assign mem_48_6_W0_en = W0_en & W0_addr_sel == 8'h30;
  assign mem_48_6_W0_mask = W0_mask[6];
  assign mem_48_7_R0_addr = R0_addr[25:0];
  assign mem_48_7_R0_clk = R0_clk;
  assign mem_48_7_R0_en = R0_en & R0_addr_sel == 8'h30;
  assign mem_48_7_W0_addr = W0_addr[25:0];
  assign mem_48_7_W0_clk = W0_clk;
  assign mem_48_7_W0_data = W0_data[63:56];
  assign mem_48_7_W0_en = W0_en & W0_addr_sel == 8'h30;
  assign mem_48_7_W0_mask = W0_mask[7];
  assign mem_49_0_R0_addr = R0_addr[25:0];
  assign mem_49_0_R0_clk = R0_clk;
  assign mem_49_0_R0_en = R0_en & R0_addr_sel == 8'h31;
  assign mem_49_0_W0_addr = W0_addr[25:0];
  assign mem_49_0_W0_clk = W0_clk;
  assign mem_49_0_W0_data = W0_data[7:0];
  assign mem_49_0_W0_en = W0_en & W0_addr_sel == 8'h31;
  assign mem_49_0_W0_mask = W0_mask[0];
  assign mem_49_1_R0_addr = R0_addr[25:0];
  assign mem_49_1_R0_clk = R0_clk;
  assign mem_49_1_R0_en = R0_en & R0_addr_sel == 8'h31;
  assign mem_49_1_W0_addr = W0_addr[25:0];
  assign mem_49_1_W0_clk = W0_clk;
  assign mem_49_1_W0_data = W0_data[15:8];
  assign mem_49_1_W0_en = W0_en & W0_addr_sel == 8'h31;
  assign mem_49_1_W0_mask = W0_mask[1];
  assign mem_49_2_R0_addr = R0_addr[25:0];
  assign mem_49_2_R0_clk = R0_clk;
  assign mem_49_2_R0_en = R0_en & R0_addr_sel == 8'h31;
  assign mem_49_2_W0_addr = W0_addr[25:0];
  assign mem_49_2_W0_clk = W0_clk;
  assign mem_49_2_W0_data = W0_data[23:16];
  assign mem_49_2_W0_en = W0_en & W0_addr_sel == 8'h31;
  assign mem_49_2_W0_mask = W0_mask[2];
  assign mem_49_3_R0_addr = R0_addr[25:0];
  assign mem_49_3_R0_clk = R0_clk;
  assign mem_49_3_R0_en = R0_en & R0_addr_sel == 8'h31;
  assign mem_49_3_W0_addr = W0_addr[25:0];
  assign mem_49_3_W0_clk = W0_clk;
  assign mem_49_3_W0_data = W0_data[31:24];
  assign mem_49_3_W0_en = W0_en & W0_addr_sel == 8'h31;
  assign mem_49_3_W0_mask = W0_mask[3];
  assign mem_49_4_R0_addr = R0_addr[25:0];
  assign mem_49_4_R0_clk = R0_clk;
  assign mem_49_4_R0_en = R0_en & R0_addr_sel == 8'h31;
  assign mem_49_4_W0_addr = W0_addr[25:0];
  assign mem_49_4_W0_clk = W0_clk;
  assign mem_49_4_W0_data = W0_data[39:32];
  assign mem_49_4_W0_en = W0_en & W0_addr_sel == 8'h31;
  assign mem_49_4_W0_mask = W0_mask[4];
  assign mem_49_5_R0_addr = R0_addr[25:0];
  assign mem_49_5_R0_clk = R0_clk;
  assign mem_49_5_R0_en = R0_en & R0_addr_sel == 8'h31;
  assign mem_49_5_W0_addr = W0_addr[25:0];
  assign mem_49_5_W0_clk = W0_clk;
  assign mem_49_5_W0_data = W0_data[47:40];
  assign mem_49_5_W0_en = W0_en & W0_addr_sel == 8'h31;
  assign mem_49_5_W0_mask = W0_mask[5];
  assign mem_49_6_R0_addr = R0_addr[25:0];
  assign mem_49_6_R0_clk = R0_clk;
  assign mem_49_6_R0_en = R0_en & R0_addr_sel == 8'h31;
  assign mem_49_6_W0_addr = W0_addr[25:0];
  assign mem_49_6_W0_clk = W0_clk;
  assign mem_49_6_W0_data = W0_data[55:48];
  assign mem_49_6_W0_en = W0_en & W0_addr_sel == 8'h31;
  assign mem_49_6_W0_mask = W0_mask[6];
  assign mem_49_7_R0_addr = R0_addr[25:0];
  assign mem_49_7_R0_clk = R0_clk;
  assign mem_49_7_R0_en = R0_en & R0_addr_sel == 8'h31;
  assign mem_49_7_W0_addr = W0_addr[25:0];
  assign mem_49_7_W0_clk = W0_clk;
  assign mem_49_7_W0_data = W0_data[63:56];
  assign mem_49_7_W0_en = W0_en & W0_addr_sel == 8'h31;
  assign mem_49_7_W0_mask = W0_mask[7];
  assign mem_50_0_R0_addr = R0_addr[25:0];
  assign mem_50_0_R0_clk = R0_clk;
  assign mem_50_0_R0_en = R0_en & R0_addr_sel == 8'h32;
  assign mem_50_0_W0_addr = W0_addr[25:0];
  assign mem_50_0_W0_clk = W0_clk;
  assign mem_50_0_W0_data = W0_data[7:0];
  assign mem_50_0_W0_en = W0_en & W0_addr_sel == 8'h32;
  assign mem_50_0_W0_mask = W0_mask[0];
  assign mem_50_1_R0_addr = R0_addr[25:0];
  assign mem_50_1_R0_clk = R0_clk;
  assign mem_50_1_R0_en = R0_en & R0_addr_sel == 8'h32;
  assign mem_50_1_W0_addr = W0_addr[25:0];
  assign mem_50_1_W0_clk = W0_clk;
  assign mem_50_1_W0_data = W0_data[15:8];
  assign mem_50_1_W0_en = W0_en & W0_addr_sel == 8'h32;
  assign mem_50_1_W0_mask = W0_mask[1];
  assign mem_50_2_R0_addr = R0_addr[25:0];
  assign mem_50_2_R0_clk = R0_clk;
  assign mem_50_2_R0_en = R0_en & R0_addr_sel == 8'h32;
  assign mem_50_2_W0_addr = W0_addr[25:0];
  assign mem_50_2_W0_clk = W0_clk;
  assign mem_50_2_W0_data = W0_data[23:16];
  assign mem_50_2_W0_en = W0_en & W0_addr_sel == 8'h32;
  assign mem_50_2_W0_mask = W0_mask[2];
  assign mem_50_3_R0_addr = R0_addr[25:0];
  assign mem_50_3_R0_clk = R0_clk;
  assign mem_50_3_R0_en = R0_en & R0_addr_sel == 8'h32;
  assign mem_50_3_W0_addr = W0_addr[25:0];
  assign mem_50_3_W0_clk = W0_clk;
  assign mem_50_3_W0_data = W0_data[31:24];
  assign mem_50_3_W0_en = W0_en & W0_addr_sel == 8'h32;
  assign mem_50_3_W0_mask = W0_mask[3];
  assign mem_50_4_R0_addr = R0_addr[25:0];
  assign mem_50_4_R0_clk = R0_clk;
  assign mem_50_4_R0_en = R0_en & R0_addr_sel == 8'h32;
  assign mem_50_4_W0_addr = W0_addr[25:0];
  assign mem_50_4_W0_clk = W0_clk;
  assign mem_50_4_W0_data = W0_data[39:32];
  assign mem_50_4_W0_en = W0_en & W0_addr_sel == 8'h32;
  assign mem_50_4_W0_mask = W0_mask[4];
  assign mem_50_5_R0_addr = R0_addr[25:0];
  assign mem_50_5_R0_clk = R0_clk;
  assign mem_50_5_R0_en = R0_en & R0_addr_sel == 8'h32;
  assign mem_50_5_W0_addr = W0_addr[25:0];
  assign mem_50_5_W0_clk = W0_clk;
  assign mem_50_5_W0_data = W0_data[47:40];
  assign mem_50_5_W0_en = W0_en & W0_addr_sel == 8'h32;
  assign mem_50_5_W0_mask = W0_mask[5];
  assign mem_50_6_R0_addr = R0_addr[25:0];
  assign mem_50_6_R0_clk = R0_clk;
  assign mem_50_6_R0_en = R0_en & R0_addr_sel == 8'h32;
  assign mem_50_6_W0_addr = W0_addr[25:0];
  assign mem_50_6_W0_clk = W0_clk;
  assign mem_50_6_W0_data = W0_data[55:48];
  assign mem_50_6_W0_en = W0_en & W0_addr_sel == 8'h32;
  assign mem_50_6_W0_mask = W0_mask[6];
  assign mem_50_7_R0_addr = R0_addr[25:0];
  assign mem_50_7_R0_clk = R0_clk;
  assign mem_50_7_R0_en = R0_en & R0_addr_sel == 8'h32;
  assign mem_50_7_W0_addr = W0_addr[25:0];
  assign mem_50_7_W0_clk = W0_clk;
  assign mem_50_7_W0_data = W0_data[63:56];
  assign mem_50_7_W0_en = W0_en & W0_addr_sel == 8'h32;
  assign mem_50_7_W0_mask = W0_mask[7];
  assign mem_51_0_R0_addr = R0_addr[25:0];
  assign mem_51_0_R0_clk = R0_clk;
  assign mem_51_0_R0_en = R0_en & R0_addr_sel == 8'h33;
  assign mem_51_0_W0_addr = W0_addr[25:0];
  assign mem_51_0_W0_clk = W0_clk;
  assign mem_51_0_W0_data = W0_data[7:0];
  assign mem_51_0_W0_en = W0_en & W0_addr_sel == 8'h33;
  assign mem_51_0_W0_mask = W0_mask[0];
  assign mem_51_1_R0_addr = R0_addr[25:0];
  assign mem_51_1_R0_clk = R0_clk;
  assign mem_51_1_R0_en = R0_en & R0_addr_sel == 8'h33;
  assign mem_51_1_W0_addr = W0_addr[25:0];
  assign mem_51_1_W0_clk = W0_clk;
  assign mem_51_1_W0_data = W0_data[15:8];
  assign mem_51_1_W0_en = W0_en & W0_addr_sel == 8'h33;
  assign mem_51_1_W0_mask = W0_mask[1];
  assign mem_51_2_R0_addr = R0_addr[25:0];
  assign mem_51_2_R0_clk = R0_clk;
  assign mem_51_2_R0_en = R0_en & R0_addr_sel == 8'h33;
  assign mem_51_2_W0_addr = W0_addr[25:0];
  assign mem_51_2_W0_clk = W0_clk;
  assign mem_51_2_W0_data = W0_data[23:16];
  assign mem_51_2_W0_en = W0_en & W0_addr_sel == 8'h33;
  assign mem_51_2_W0_mask = W0_mask[2];
  assign mem_51_3_R0_addr = R0_addr[25:0];
  assign mem_51_3_R0_clk = R0_clk;
  assign mem_51_3_R0_en = R0_en & R0_addr_sel == 8'h33;
  assign mem_51_3_W0_addr = W0_addr[25:0];
  assign mem_51_3_W0_clk = W0_clk;
  assign mem_51_3_W0_data = W0_data[31:24];
  assign mem_51_3_W0_en = W0_en & W0_addr_sel == 8'h33;
  assign mem_51_3_W0_mask = W0_mask[3];
  assign mem_51_4_R0_addr = R0_addr[25:0];
  assign mem_51_4_R0_clk = R0_clk;
  assign mem_51_4_R0_en = R0_en & R0_addr_sel == 8'h33;
  assign mem_51_4_W0_addr = W0_addr[25:0];
  assign mem_51_4_W0_clk = W0_clk;
  assign mem_51_4_W0_data = W0_data[39:32];
  assign mem_51_4_W0_en = W0_en & W0_addr_sel == 8'h33;
  assign mem_51_4_W0_mask = W0_mask[4];
  assign mem_51_5_R0_addr = R0_addr[25:0];
  assign mem_51_5_R0_clk = R0_clk;
  assign mem_51_5_R0_en = R0_en & R0_addr_sel == 8'h33;
  assign mem_51_5_W0_addr = W0_addr[25:0];
  assign mem_51_5_W0_clk = W0_clk;
  assign mem_51_5_W0_data = W0_data[47:40];
  assign mem_51_5_W0_en = W0_en & W0_addr_sel == 8'h33;
  assign mem_51_5_W0_mask = W0_mask[5];
  assign mem_51_6_R0_addr = R0_addr[25:0];
  assign mem_51_6_R0_clk = R0_clk;
  assign mem_51_6_R0_en = R0_en & R0_addr_sel == 8'h33;
  assign mem_51_6_W0_addr = W0_addr[25:0];
  assign mem_51_6_W0_clk = W0_clk;
  assign mem_51_6_W0_data = W0_data[55:48];
  assign mem_51_6_W0_en = W0_en & W0_addr_sel == 8'h33;
  assign mem_51_6_W0_mask = W0_mask[6];
  assign mem_51_7_R0_addr = R0_addr[25:0];
  assign mem_51_7_R0_clk = R0_clk;
  assign mem_51_7_R0_en = R0_en & R0_addr_sel == 8'h33;
  assign mem_51_7_W0_addr = W0_addr[25:0];
  assign mem_51_7_W0_clk = W0_clk;
  assign mem_51_7_W0_data = W0_data[63:56];
  assign mem_51_7_W0_en = W0_en & W0_addr_sel == 8'h33;
  assign mem_51_7_W0_mask = W0_mask[7];
  assign mem_52_0_R0_addr = R0_addr[25:0];
  assign mem_52_0_R0_clk = R0_clk;
  assign mem_52_0_R0_en = R0_en & R0_addr_sel == 8'h34;
  assign mem_52_0_W0_addr = W0_addr[25:0];
  assign mem_52_0_W0_clk = W0_clk;
  assign mem_52_0_W0_data = W0_data[7:0];
  assign mem_52_0_W0_en = W0_en & W0_addr_sel == 8'h34;
  assign mem_52_0_W0_mask = W0_mask[0];
  assign mem_52_1_R0_addr = R0_addr[25:0];
  assign mem_52_1_R0_clk = R0_clk;
  assign mem_52_1_R0_en = R0_en & R0_addr_sel == 8'h34;
  assign mem_52_1_W0_addr = W0_addr[25:0];
  assign mem_52_1_W0_clk = W0_clk;
  assign mem_52_1_W0_data = W0_data[15:8];
  assign mem_52_1_W0_en = W0_en & W0_addr_sel == 8'h34;
  assign mem_52_1_W0_mask = W0_mask[1];
  assign mem_52_2_R0_addr = R0_addr[25:0];
  assign mem_52_2_R0_clk = R0_clk;
  assign mem_52_2_R0_en = R0_en & R0_addr_sel == 8'h34;
  assign mem_52_2_W0_addr = W0_addr[25:0];
  assign mem_52_2_W0_clk = W0_clk;
  assign mem_52_2_W0_data = W0_data[23:16];
  assign mem_52_2_W0_en = W0_en & W0_addr_sel == 8'h34;
  assign mem_52_2_W0_mask = W0_mask[2];
  assign mem_52_3_R0_addr = R0_addr[25:0];
  assign mem_52_3_R0_clk = R0_clk;
  assign mem_52_3_R0_en = R0_en & R0_addr_sel == 8'h34;
  assign mem_52_3_W0_addr = W0_addr[25:0];
  assign mem_52_3_W0_clk = W0_clk;
  assign mem_52_3_W0_data = W0_data[31:24];
  assign mem_52_3_W0_en = W0_en & W0_addr_sel == 8'h34;
  assign mem_52_3_W0_mask = W0_mask[3];
  assign mem_52_4_R0_addr = R0_addr[25:0];
  assign mem_52_4_R0_clk = R0_clk;
  assign mem_52_4_R0_en = R0_en & R0_addr_sel == 8'h34;
  assign mem_52_4_W0_addr = W0_addr[25:0];
  assign mem_52_4_W0_clk = W0_clk;
  assign mem_52_4_W0_data = W0_data[39:32];
  assign mem_52_4_W0_en = W0_en & W0_addr_sel == 8'h34;
  assign mem_52_4_W0_mask = W0_mask[4];
  assign mem_52_5_R0_addr = R0_addr[25:0];
  assign mem_52_5_R0_clk = R0_clk;
  assign mem_52_5_R0_en = R0_en & R0_addr_sel == 8'h34;
  assign mem_52_5_W0_addr = W0_addr[25:0];
  assign mem_52_5_W0_clk = W0_clk;
  assign mem_52_5_W0_data = W0_data[47:40];
  assign mem_52_5_W0_en = W0_en & W0_addr_sel == 8'h34;
  assign mem_52_5_W0_mask = W0_mask[5];
  assign mem_52_6_R0_addr = R0_addr[25:0];
  assign mem_52_6_R0_clk = R0_clk;
  assign mem_52_6_R0_en = R0_en & R0_addr_sel == 8'h34;
  assign mem_52_6_W0_addr = W0_addr[25:0];
  assign mem_52_6_W0_clk = W0_clk;
  assign mem_52_6_W0_data = W0_data[55:48];
  assign mem_52_6_W0_en = W0_en & W0_addr_sel == 8'h34;
  assign mem_52_6_W0_mask = W0_mask[6];
  assign mem_52_7_R0_addr = R0_addr[25:0];
  assign mem_52_7_R0_clk = R0_clk;
  assign mem_52_7_R0_en = R0_en & R0_addr_sel == 8'h34;
  assign mem_52_7_W0_addr = W0_addr[25:0];
  assign mem_52_7_W0_clk = W0_clk;
  assign mem_52_7_W0_data = W0_data[63:56];
  assign mem_52_7_W0_en = W0_en & W0_addr_sel == 8'h34;
  assign mem_52_7_W0_mask = W0_mask[7];
  assign mem_53_0_R0_addr = R0_addr[25:0];
  assign mem_53_0_R0_clk = R0_clk;
  assign mem_53_0_R0_en = R0_en & R0_addr_sel == 8'h35;
  assign mem_53_0_W0_addr = W0_addr[25:0];
  assign mem_53_0_W0_clk = W0_clk;
  assign mem_53_0_W0_data = W0_data[7:0];
  assign mem_53_0_W0_en = W0_en & W0_addr_sel == 8'h35;
  assign mem_53_0_W0_mask = W0_mask[0];
  assign mem_53_1_R0_addr = R0_addr[25:0];
  assign mem_53_1_R0_clk = R0_clk;
  assign mem_53_1_R0_en = R0_en & R0_addr_sel == 8'h35;
  assign mem_53_1_W0_addr = W0_addr[25:0];
  assign mem_53_1_W0_clk = W0_clk;
  assign mem_53_1_W0_data = W0_data[15:8];
  assign mem_53_1_W0_en = W0_en & W0_addr_sel == 8'h35;
  assign mem_53_1_W0_mask = W0_mask[1];
  assign mem_53_2_R0_addr = R0_addr[25:0];
  assign mem_53_2_R0_clk = R0_clk;
  assign mem_53_2_R0_en = R0_en & R0_addr_sel == 8'h35;
  assign mem_53_2_W0_addr = W0_addr[25:0];
  assign mem_53_2_W0_clk = W0_clk;
  assign mem_53_2_W0_data = W0_data[23:16];
  assign mem_53_2_W0_en = W0_en & W0_addr_sel == 8'h35;
  assign mem_53_2_W0_mask = W0_mask[2];
  assign mem_53_3_R0_addr = R0_addr[25:0];
  assign mem_53_3_R0_clk = R0_clk;
  assign mem_53_3_R0_en = R0_en & R0_addr_sel == 8'h35;
  assign mem_53_3_W0_addr = W0_addr[25:0];
  assign mem_53_3_W0_clk = W0_clk;
  assign mem_53_3_W0_data = W0_data[31:24];
  assign mem_53_3_W0_en = W0_en & W0_addr_sel == 8'h35;
  assign mem_53_3_W0_mask = W0_mask[3];
  assign mem_53_4_R0_addr = R0_addr[25:0];
  assign mem_53_4_R0_clk = R0_clk;
  assign mem_53_4_R0_en = R0_en & R0_addr_sel == 8'h35;
  assign mem_53_4_W0_addr = W0_addr[25:0];
  assign mem_53_4_W0_clk = W0_clk;
  assign mem_53_4_W0_data = W0_data[39:32];
  assign mem_53_4_W0_en = W0_en & W0_addr_sel == 8'h35;
  assign mem_53_4_W0_mask = W0_mask[4];
  assign mem_53_5_R0_addr = R0_addr[25:0];
  assign mem_53_5_R0_clk = R0_clk;
  assign mem_53_5_R0_en = R0_en & R0_addr_sel == 8'h35;
  assign mem_53_5_W0_addr = W0_addr[25:0];
  assign mem_53_5_W0_clk = W0_clk;
  assign mem_53_5_W0_data = W0_data[47:40];
  assign mem_53_5_W0_en = W0_en & W0_addr_sel == 8'h35;
  assign mem_53_5_W0_mask = W0_mask[5];
  assign mem_53_6_R0_addr = R0_addr[25:0];
  assign mem_53_6_R0_clk = R0_clk;
  assign mem_53_6_R0_en = R0_en & R0_addr_sel == 8'h35;
  assign mem_53_6_W0_addr = W0_addr[25:0];
  assign mem_53_6_W0_clk = W0_clk;
  assign mem_53_6_W0_data = W0_data[55:48];
  assign mem_53_6_W0_en = W0_en & W0_addr_sel == 8'h35;
  assign mem_53_6_W0_mask = W0_mask[6];
  assign mem_53_7_R0_addr = R0_addr[25:0];
  assign mem_53_7_R0_clk = R0_clk;
  assign mem_53_7_R0_en = R0_en & R0_addr_sel == 8'h35;
  assign mem_53_7_W0_addr = W0_addr[25:0];
  assign mem_53_7_W0_clk = W0_clk;
  assign mem_53_7_W0_data = W0_data[63:56];
  assign mem_53_7_W0_en = W0_en & W0_addr_sel == 8'h35;
  assign mem_53_7_W0_mask = W0_mask[7];
  assign mem_54_0_R0_addr = R0_addr[25:0];
  assign mem_54_0_R0_clk = R0_clk;
  assign mem_54_0_R0_en = R0_en & R0_addr_sel == 8'h36;
  assign mem_54_0_W0_addr = W0_addr[25:0];
  assign mem_54_0_W0_clk = W0_clk;
  assign mem_54_0_W0_data = W0_data[7:0];
  assign mem_54_0_W0_en = W0_en & W0_addr_sel == 8'h36;
  assign mem_54_0_W0_mask = W0_mask[0];
  assign mem_54_1_R0_addr = R0_addr[25:0];
  assign mem_54_1_R0_clk = R0_clk;
  assign mem_54_1_R0_en = R0_en & R0_addr_sel == 8'h36;
  assign mem_54_1_W0_addr = W0_addr[25:0];
  assign mem_54_1_W0_clk = W0_clk;
  assign mem_54_1_W0_data = W0_data[15:8];
  assign mem_54_1_W0_en = W0_en & W0_addr_sel == 8'h36;
  assign mem_54_1_W0_mask = W0_mask[1];
  assign mem_54_2_R0_addr = R0_addr[25:0];
  assign mem_54_2_R0_clk = R0_clk;
  assign mem_54_2_R0_en = R0_en & R0_addr_sel == 8'h36;
  assign mem_54_2_W0_addr = W0_addr[25:0];
  assign mem_54_2_W0_clk = W0_clk;
  assign mem_54_2_W0_data = W0_data[23:16];
  assign mem_54_2_W0_en = W0_en & W0_addr_sel == 8'h36;
  assign mem_54_2_W0_mask = W0_mask[2];
  assign mem_54_3_R0_addr = R0_addr[25:0];
  assign mem_54_3_R0_clk = R0_clk;
  assign mem_54_3_R0_en = R0_en & R0_addr_sel == 8'h36;
  assign mem_54_3_W0_addr = W0_addr[25:0];
  assign mem_54_3_W0_clk = W0_clk;
  assign mem_54_3_W0_data = W0_data[31:24];
  assign mem_54_3_W0_en = W0_en & W0_addr_sel == 8'h36;
  assign mem_54_3_W0_mask = W0_mask[3];
  assign mem_54_4_R0_addr = R0_addr[25:0];
  assign mem_54_4_R0_clk = R0_clk;
  assign mem_54_4_R0_en = R0_en & R0_addr_sel == 8'h36;
  assign mem_54_4_W0_addr = W0_addr[25:0];
  assign mem_54_4_W0_clk = W0_clk;
  assign mem_54_4_W0_data = W0_data[39:32];
  assign mem_54_4_W0_en = W0_en & W0_addr_sel == 8'h36;
  assign mem_54_4_W0_mask = W0_mask[4];
  assign mem_54_5_R0_addr = R0_addr[25:0];
  assign mem_54_5_R0_clk = R0_clk;
  assign mem_54_5_R0_en = R0_en & R0_addr_sel == 8'h36;
  assign mem_54_5_W0_addr = W0_addr[25:0];
  assign mem_54_5_W0_clk = W0_clk;
  assign mem_54_5_W0_data = W0_data[47:40];
  assign mem_54_5_W0_en = W0_en & W0_addr_sel == 8'h36;
  assign mem_54_5_W0_mask = W0_mask[5];
  assign mem_54_6_R0_addr = R0_addr[25:0];
  assign mem_54_6_R0_clk = R0_clk;
  assign mem_54_6_R0_en = R0_en & R0_addr_sel == 8'h36;
  assign mem_54_6_W0_addr = W0_addr[25:0];
  assign mem_54_6_W0_clk = W0_clk;
  assign mem_54_6_W0_data = W0_data[55:48];
  assign mem_54_6_W0_en = W0_en & W0_addr_sel == 8'h36;
  assign mem_54_6_W0_mask = W0_mask[6];
  assign mem_54_7_R0_addr = R0_addr[25:0];
  assign mem_54_7_R0_clk = R0_clk;
  assign mem_54_7_R0_en = R0_en & R0_addr_sel == 8'h36;
  assign mem_54_7_W0_addr = W0_addr[25:0];
  assign mem_54_7_W0_clk = W0_clk;
  assign mem_54_7_W0_data = W0_data[63:56];
  assign mem_54_7_W0_en = W0_en & W0_addr_sel == 8'h36;
  assign mem_54_7_W0_mask = W0_mask[7];
  assign mem_55_0_R0_addr = R0_addr[25:0];
  assign mem_55_0_R0_clk = R0_clk;
  assign mem_55_0_R0_en = R0_en & R0_addr_sel == 8'h37;
  assign mem_55_0_W0_addr = W0_addr[25:0];
  assign mem_55_0_W0_clk = W0_clk;
  assign mem_55_0_W0_data = W0_data[7:0];
  assign mem_55_0_W0_en = W0_en & W0_addr_sel == 8'h37;
  assign mem_55_0_W0_mask = W0_mask[0];
  assign mem_55_1_R0_addr = R0_addr[25:0];
  assign mem_55_1_R0_clk = R0_clk;
  assign mem_55_1_R0_en = R0_en & R0_addr_sel == 8'h37;
  assign mem_55_1_W0_addr = W0_addr[25:0];
  assign mem_55_1_W0_clk = W0_clk;
  assign mem_55_1_W0_data = W0_data[15:8];
  assign mem_55_1_W0_en = W0_en & W0_addr_sel == 8'h37;
  assign mem_55_1_W0_mask = W0_mask[1];
  assign mem_55_2_R0_addr = R0_addr[25:0];
  assign mem_55_2_R0_clk = R0_clk;
  assign mem_55_2_R0_en = R0_en & R0_addr_sel == 8'h37;
  assign mem_55_2_W0_addr = W0_addr[25:0];
  assign mem_55_2_W0_clk = W0_clk;
  assign mem_55_2_W0_data = W0_data[23:16];
  assign mem_55_2_W0_en = W0_en & W0_addr_sel == 8'h37;
  assign mem_55_2_W0_mask = W0_mask[2];
  assign mem_55_3_R0_addr = R0_addr[25:0];
  assign mem_55_3_R0_clk = R0_clk;
  assign mem_55_3_R0_en = R0_en & R0_addr_sel == 8'h37;
  assign mem_55_3_W0_addr = W0_addr[25:0];
  assign mem_55_3_W0_clk = W0_clk;
  assign mem_55_3_W0_data = W0_data[31:24];
  assign mem_55_3_W0_en = W0_en & W0_addr_sel == 8'h37;
  assign mem_55_3_W0_mask = W0_mask[3];
  assign mem_55_4_R0_addr = R0_addr[25:0];
  assign mem_55_4_R0_clk = R0_clk;
  assign mem_55_4_R0_en = R0_en & R0_addr_sel == 8'h37;
  assign mem_55_4_W0_addr = W0_addr[25:0];
  assign mem_55_4_W0_clk = W0_clk;
  assign mem_55_4_W0_data = W0_data[39:32];
  assign mem_55_4_W0_en = W0_en & W0_addr_sel == 8'h37;
  assign mem_55_4_W0_mask = W0_mask[4];
  assign mem_55_5_R0_addr = R0_addr[25:0];
  assign mem_55_5_R0_clk = R0_clk;
  assign mem_55_5_R0_en = R0_en & R0_addr_sel == 8'h37;
  assign mem_55_5_W0_addr = W0_addr[25:0];
  assign mem_55_5_W0_clk = W0_clk;
  assign mem_55_5_W0_data = W0_data[47:40];
  assign mem_55_5_W0_en = W0_en & W0_addr_sel == 8'h37;
  assign mem_55_5_W0_mask = W0_mask[5];
  assign mem_55_6_R0_addr = R0_addr[25:0];
  assign mem_55_6_R0_clk = R0_clk;
  assign mem_55_6_R0_en = R0_en & R0_addr_sel == 8'h37;
  assign mem_55_6_W0_addr = W0_addr[25:0];
  assign mem_55_6_W0_clk = W0_clk;
  assign mem_55_6_W0_data = W0_data[55:48];
  assign mem_55_6_W0_en = W0_en & W0_addr_sel == 8'h37;
  assign mem_55_6_W0_mask = W0_mask[6];
  assign mem_55_7_R0_addr = R0_addr[25:0];
  assign mem_55_7_R0_clk = R0_clk;
  assign mem_55_7_R0_en = R0_en & R0_addr_sel == 8'h37;
  assign mem_55_7_W0_addr = W0_addr[25:0];
  assign mem_55_7_W0_clk = W0_clk;
  assign mem_55_7_W0_data = W0_data[63:56];
  assign mem_55_7_W0_en = W0_en & W0_addr_sel == 8'h37;
  assign mem_55_7_W0_mask = W0_mask[7];
  assign mem_56_0_R0_addr = R0_addr[25:0];
  assign mem_56_0_R0_clk = R0_clk;
  assign mem_56_0_R0_en = R0_en & R0_addr_sel == 8'h38;
  assign mem_56_0_W0_addr = W0_addr[25:0];
  assign mem_56_0_W0_clk = W0_clk;
  assign mem_56_0_W0_data = W0_data[7:0];
  assign mem_56_0_W0_en = W0_en & W0_addr_sel == 8'h38;
  assign mem_56_0_W0_mask = W0_mask[0];
  assign mem_56_1_R0_addr = R0_addr[25:0];
  assign mem_56_1_R0_clk = R0_clk;
  assign mem_56_1_R0_en = R0_en & R0_addr_sel == 8'h38;
  assign mem_56_1_W0_addr = W0_addr[25:0];
  assign mem_56_1_W0_clk = W0_clk;
  assign mem_56_1_W0_data = W0_data[15:8];
  assign mem_56_1_W0_en = W0_en & W0_addr_sel == 8'h38;
  assign mem_56_1_W0_mask = W0_mask[1];
  assign mem_56_2_R0_addr = R0_addr[25:0];
  assign mem_56_2_R0_clk = R0_clk;
  assign mem_56_2_R0_en = R0_en & R0_addr_sel == 8'h38;
  assign mem_56_2_W0_addr = W0_addr[25:0];
  assign mem_56_2_W0_clk = W0_clk;
  assign mem_56_2_W0_data = W0_data[23:16];
  assign mem_56_2_W0_en = W0_en & W0_addr_sel == 8'h38;
  assign mem_56_2_W0_mask = W0_mask[2];
  assign mem_56_3_R0_addr = R0_addr[25:0];
  assign mem_56_3_R0_clk = R0_clk;
  assign mem_56_3_R0_en = R0_en & R0_addr_sel == 8'h38;
  assign mem_56_3_W0_addr = W0_addr[25:0];
  assign mem_56_3_W0_clk = W0_clk;
  assign mem_56_3_W0_data = W0_data[31:24];
  assign mem_56_3_W0_en = W0_en & W0_addr_sel == 8'h38;
  assign mem_56_3_W0_mask = W0_mask[3];
  assign mem_56_4_R0_addr = R0_addr[25:0];
  assign mem_56_4_R0_clk = R0_clk;
  assign mem_56_4_R0_en = R0_en & R0_addr_sel == 8'h38;
  assign mem_56_4_W0_addr = W0_addr[25:0];
  assign mem_56_4_W0_clk = W0_clk;
  assign mem_56_4_W0_data = W0_data[39:32];
  assign mem_56_4_W0_en = W0_en & W0_addr_sel == 8'h38;
  assign mem_56_4_W0_mask = W0_mask[4];
  assign mem_56_5_R0_addr = R0_addr[25:0];
  assign mem_56_5_R0_clk = R0_clk;
  assign mem_56_5_R0_en = R0_en & R0_addr_sel == 8'h38;
  assign mem_56_5_W0_addr = W0_addr[25:0];
  assign mem_56_5_W0_clk = W0_clk;
  assign mem_56_5_W0_data = W0_data[47:40];
  assign mem_56_5_W0_en = W0_en & W0_addr_sel == 8'h38;
  assign mem_56_5_W0_mask = W0_mask[5];
  assign mem_56_6_R0_addr = R0_addr[25:0];
  assign mem_56_6_R0_clk = R0_clk;
  assign mem_56_6_R0_en = R0_en & R0_addr_sel == 8'h38;
  assign mem_56_6_W0_addr = W0_addr[25:0];
  assign mem_56_6_W0_clk = W0_clk;
  assign mem_56_6_W0_data = W0_data[55:48];
  assign mem_56_6_W0_en = W0_en & W0_addr_sel == 8'h38;
  assign mem_56_6_W0_mask = W0_mask[6];
  assign mem_56_7_R0_addr = R0_addr[25:0];
  assign mem_56_7_R0_clk = R0_clk;
  assign mem_56_7_R0_en = R0_en & R0_addr_sel == 8'h38;
  assign mem_56_7_W0_addr = W0_addr[25:0];
  assign mem_56_7_W0_clk = W0_clk;
  assign mem_56_7_W0_data = W0_data[63:56];
  assign mem_56_7_W0_en = W0_en & W0_addr_sel == 8'h38;
  assign mem_56_7_W0_mask = W0_mask[7];
  assign mem_57_0_R0_addr = R0_addr[25:0];
  assign mem_57_0_R0_clk = R0_clk;
  assign mem_57_0_R0_en = R0_en & R0_addr_sel == 8'h39;
  assign mem_57_0_W0_addr = W0_addr[25:0];
  assign mem_57_0_W0_clk = W0_clk;
  assign mem_57_0_W0_data = W0_data[7:0];
  assign mem_57_0_W0_en = W0_en & W0_addr_sel == 8'h39;
  assign mem_57_0_W0_mask = W0_mask[0];
  assign mem_57_1_R0_addr = R0_addr[25:0];
  assign mem_57_1_R0_clk = R0_clk;
  assign mem_57_1_R0_en = R0_en & R0_addr_sel == 8'h39;
  assign mem_57_1_W0_addr = W0_addr[25:0];
  assign mem_57_1_W0_clk = W0_clk;
  assign mem_57_1_W0_data = W0_data[15:8];
  assign mem_57_1_W0_en = W0_en & W0_addr_sel == 8'h39;
  assign mem_57_1_W0_mask = W0_mask[1];
  assign mem_57_2_R0_addr = R0_addr[25:0];
  assign mem_57_2_R0_clk = R0_clk;
  assign mem_57_2_R0_en = R0_en & R0_addr_sel == 8'h39;
  assign mem_57_2_W0_addr = W0_addr[25:0];
  assign mem_57_2_W0_clk = W0_clk;
  assign mem_57_2_W0_data = W0_data[23:16];
  assign mem_57_2_W0_en = W0_en & W0_addr_sel == 8'h39;
  assign mem_57_2_W0_mask = W0_mask[2];
  assign mem_57_3_R0_addr = R0_addr[25:0];
  assign mem_57_3_R0_clk = R0_clk;
  assign mem_57_3_R0_en = R0_en & R0_addr_sel == 8'h39;
  assign mem_57_3_W0_addr = W0_addr[25:0];
  assign mem_57_3_W0_clk = W0_clk;
  assign mem_57_3_W0_data = W0_data[31:24];
  assign mem_57_3_W0_en = W0_en & W0_addr_sel == 8'h39;
  assign mem_57_3_W0_mask = W0_mask[3];
  assign mem_57_4_R0_addr = R0_addr[25:0];
  assign mem_57_4_R0_clk = R0_clk;
  assign mem_57_4_R0_en = R0_en & R0_addr_sel == 8'h39;
  assign mem_57_4_W0_addr = W0_addr[25:0];
  assign mem_57_4_W0_clk = W0_clk;
  assign mem_57_4_W0_data = W0_data[39:32];
  assign mem_57_4_W0_en = W0_en & W0_addr_sel == 8'h39;
  assign mem_57_4_W0_mask = W0_mask[4];
  assign mem_57_5_R0_addr = R0_addr[25:0];
  assign mem_57_5_R0_clk = R0_clk;
  assign mem_57_5_R0_en = R0_en & R0_addr_sel == 8'h39;
  assign mem_57_5_W0_addr = W0_addr[25:0];
  assign mem_57_5_W0_clk = W0_clk;
  assign mem_57_5_W0_data = W0_data[47:40];
  assign mem_57_5_W0_en = W0_en & W0_addr_sel == 8'h39;
  assign mem_57_5_W0_mask = W0_mask[5];
  assign mem_57_6_R0_addr = R0_addr[25:0];
  assign mem_57_6_R0_clk = R0_clk;
  assign mem_57_6_R0_en = R0_en & R0_addr_sel == 8'h39;
  assign mem_57_6_W0_addr = W0_addr[25:0];
  assign mem_57_6_W0_clk = W0_clk;
  assign mem_57_6_W0_data = W0_data[55:48];
  assign mem_57_6_W0_en = W0_en & W0_addr_sel == 8'h39;
  assign mem_57_6_W0_mask = W0_mask[6];
  assign mem_57_7_R0_addr = R0_addr[25:0];
  assign mem_57_7_R0_clk = R0_clk;
  assign mem_57_7_R0_en = R0_en & R0_addr_sel == 8'h39;
  assign mem_57_7_W0_addr = W0_addr[25:0];
  assign mem_57_7_W0_clk = W0_clk;
  assign mem_57_7_W0_data = W0_data[63:56];
  assign mem_57_7_W0_en = W0_en & W0_addr_sel == 8'h39;
  assign mem_57_7_W0_mask = W0_mask[7];
  assign mem_58_0_R0_addr = R0_addr[25:0];
  assign mem_58_0_R0_clk = R0_clk;
  assign mem_58_0_R0_en = R0_en & R0_addr_sel == 8'h3a;
  assign mem_58_0_W0_addr = W0_addr[25:0];
  assign mem_58_0_W0_clk = W0_clk;
  assign mem_58_0_W0_data = W0_data[7:0];
  assign mem_58_0_W0_en = W0_en & W0_addr_sel == 8'h3a;
  assign mem_58_0_W0_mask = W0_mask[0];
  assign mem_58_1_R0_addr = R0_addr[25:0];
  assign mem_58_1_R0_clk = R0_clk;
  assign mem_58_1_R0_en = R0_en & R0_addr_sel == 8'h3a;
  assign mem_58_1_W0_addr = W0_addr[25:0];
  assign mem_58_1_W0_clk = W0_clk;
  assign mem_58_1_W0_data = W0_data[15:8];
  assign mem_58_1_W0_en = W0_en & W0_addr_sel == 8'h3a;
  assign mem_58_1_W0_mask = W0_mask[1];
  assign mem_58_2_R0_addr = R0_addr[25:0];
  assign mem_58_2_R0_clk = R0_clk;
  assign mem_58_2_R0_en = R0_en & R0_addr_sel == 8'h3a;
  assign mem_58_2_W0_addr = W0_addr[25:0];
  assign mem_58_2_W0_clk = W0_clk;
  assign mem_58_2_W0_data = W0_data[23:16];
  assign mem_58_2_W0_en = W0_en & W0_addr_sel == 8'h3a;
  assign mem_58_2_W0_mask = W0_mask[2];
  assign mem_58_3_R0_addr = R0_addr[25:0];
  assign mem_58_3_R0_clk = R0_clk;
  assign mem_58_3_R0_en = R0_en & R0_addr_sel == 8'h3a;
  assign mem_58_3_W0_addr = W0_addr[25:0];
  assign mem_58_3_W0_clk = W0_clk;
  assign mem_58_3_W0_data = W0_data[31:24];
  assign mem_58_3_W0_en = W0_en & W0_addr_sel == 8'h3a;
  assign mem_58_3_W0_mask = W0_mask[3];
  assign mem_58_4_R0_addr = R0_addr[25:0];
  assign mem_58_4_R0_clk = R0_clk;
  assign mem_58_4_R0_en = R0_en & R0_addr_sel == 8'h3a;
  assign mem_58_4_W0_addr = W0_addr[25:0];
  assign mem_58_4_W0_clk = W0_clk;
  assign mem_58_4_W0_data = W0_data[39:32];
  assign mem_58_4_W0_en = W0_en & W0_addr_sel == 8'h3a;
  assign mem_58_4_W0_mask = W0_mask[4];
  assign mem_58_5_R0_addr = R0_addr[25:0];
  assign mem_58_5_R0_clk = R0_clk;
  assign mem_58_5_R0_en = R0_en & R0_addr_sel == 8'h3a;
  assign mem_58_5_W0_addr = W0_addr[25:0];
  assign mem_58_5_W0_clk = W0_clk;
  assign mem_58_5_W0_data = W0_data[47:40];
  assign mem_58_5_W0_en = W0_en & W0_addr_sel == 8'h3a;
  assign mem_58_5_W0_mask = W0_mask[5];
  assign mem_58_6_R0_addr = R0_addr[25:0];
  assign mem_58_6_R0_clk = R0_clk;
  assign mem_58_6_R0_en = R0_en & R0_addr_sel == 8'h3a;
  assign mem_58_6_W0_addr = W0_addr[25:0];
  assign mem_58_6_W0_clk = W0_clk;
  assign mem_58_6_W0_data = W0_data[55:48];
  assign mem_58_6_W0_en = W0_en & W0_addr_sel == 8'h3a;
  assign mem_58_6_W0_mask = W0_mask[6];
  assign mem_58_7_R0_addr = R0_addr[25:0];
  assign mem_58_7_R0_clk = R0_clk;
  assign mem_58_7_R0_en = R0_en & R0_addr_sel == 8'h3a;
  assign mem_58_7_W0_addr = W0_addr[25:0];
  assign mem_58_7_W0_clk = W0_clk;
  assign mem_58_7_W0_data = W0_data[63:56];
  assign mem_58_7_W0_en = W0_en & W0_addr_sel == 8'h3a;
  assign mem_58_7_W0_mask = W0_mask[7];
  assign mem_59_0_R0_addr = R0_addr[25:0];
  assign mem_59_0_R0_clk = R0_clk;
  assign mem_59_0_R0_en = R0_en & R0_addr_sel == 8'h3b;
  assign mem_59_0_W0_addr = W0_addr[25:0];
  assign mem_59_0_W0_clk = W0_clk;
  assign mem_59_0_W0_data = W0_data[7:0];
  assign mem_59_0_W0_en = W0_en & W0_addr_sel == 8'h3b;
  assign mem_59_0_W0_mask = W0_mask[0];
  assign mem_59_1_R0_addr = R0_addr[25:0];
  assign mem_59_1_R0_clk = R0_clk;
  assign mem_59_1_R0_en = R0_en & R0_addr_sel == 8'h3b;
  assign mem_59_1_W0_addr = W0_addr[25:0];
  assign mem_59_1_W0_clk = W0_clk;
  assign mem_59_1_W0_data = W0_data[15:8];
  assign mem_59_1_W0_en = W0_en & W0_addr_sel == 8'h3b;
  assign mem_59_1_W0_mask = W0_mask[1];
  assign mem_59_2_R0_addr = R0_addr[25:0];
  assign mem_59_2_R0_clk = R0_clk;
  assign mem_59_2_R0_en = R0_en & R0_addr_sel == 8'h3b;
  assign mem_59_2_W0_addr = W0_addr[25:0];
  assign mem_59_2_W0_clk = W0_clk;
  assign mem_59_2_W0_data = W0_data[23:16];
  assign mem_59_2_W0_en = W0_en & W0_addr_sel == 8'h3b;
  assign mem_59_2_W0_mask = W0_mask[2];
  assign mem_59_3_R0_addr = R0_addr[25:0];
  assign mem_59_3_R0_clk = R0_clk;
  assign mem_59_3_R0_en = R0_en & R0_addr_sel == 8'h3b;
  assign mem_59_3_W0_addr = W0_addr[25:0];
  assign mem_59_3_W0_clk = W0_clk;
  assign mem_59_3_W0_data = W0_data[31:24];
  assign mem_59_3_W0_en = W0_en & W0_addr_sel == 8'h3b;
  assign mem_59_3_W0_mask = W0_mask[3];
  assign mem_59_4_R0_addr = R0_addr[25:0];
  assign mem_59_4_R0_clk = R0_clk;
  assign mem_59_4_R0_en = R0_en & R0_addr_sel == 8'h3b;
  assign mem_59_4_W0_addr = W0_addr[25:0];
  assign mem_59_4_W0_clk = W0_clk;
  assign mem_59_4_W0_data = W0_data[39:32];
  assign mem_59_4_W0_en = W0_en & W0_addr_sel == 8'h3b;
  assign mem_59_4_W0_mask = W0_mask[4];
  assign mem_59_5_R0_addr = R0_addr[25:0];
  assign mem_59_5_R0_clk = R0_clk;
  assign mem_59_5_R0_en = R0_en & R0_addr_sel == 8'h3b;
  assign mem_59_5_W0_addr = W0_addr[25:0];
  assign mem_59_5_W0_clk = W0_clk;
  assign mem_59_5_W0_data = W0_data[47:40];
  assign mem_59_5_W0_en = W0_en & W0_addr_sel == 8'h3b;
  assign mem_59_5_W0_mask = W0_mask[5];
  assign mem_59_6_R0_addr = R0_addr[25:0];
  assign mem_59_6_R0_clk = R0_clk;
  assign mem_59_6_R0_en = R0_en & R0_addr_sel == 8'h3b;
  assign mem_59_6_W0_addr = W0_addr[25:0];
  assign mem_59_6_W0_clk = W0_clk;
  assign mem_59_6_W0_data = W0_data[55:48];
  assign mem_59_6_W0_en = W0_en & W0_addr_sel == 8'h3b;
  assign mem_59_6_W0_mask = W0_mask[6];
  assign mem_59_7_R0_addr = R0_addr[25:0];
  assign mem_59_7_R0_clk = R0_clk;
  assign mem_59_7_R0_en = R0_en & R0_addr_sel == 8'h3b;
  assign mem_59_7_W0_addr = W0_addr[25:0];
  assign mem_59_7_W0_clk = W0_clk;
  assign mem_59_7_W0_data = W0_data[63:56];
  assign mem_59_7_W0_en = W0_en & W0_addr_sel == 8'h3b;
  assign mem_59_7_W0_mask = W0_mask[7];
  assign mem_60_0_R0_addr = R0_addr[25:0];
  assign mem_60_0_R0_clk = R0_clk;
  assign mem_60_0_R0_en = R0_en & R0_addr_sel == 8'h3c;
  assign mem_60_0_W0_addr = W0_addr[25:0];
  assign mem_60_0_W0_clk = W0_clk;
  assign mem_60_0_W0_data = W0_data[7:0];
  assign mem_60_0_W0_en = W0_en & W0_addr_sel == 8'h3c;
  assign mem_60_0_W0_mask = W0_mask[0];
  assign mem_60_1_R0_addr = R0_addr[25:0];
  assign mem_60_1_R0_clk = R0_clk;
  assign mem_60_1_R0_en = R0_en & R0_addr_sel == 8'h3c;
  assign mem_60_1_W0_addr = W0_addr[25:0];
  assign mem_60_1_W0_clk = W0_clk;
  assign mem_60_1_W0_data = W0_data[15:8];
  assign mem_60_1_W0_en = W0_en & W0_addr_sel == 8'h3c;
  assign mem_60_1_W0_mask = W0_mask[1];
  assign mem_60_2_R0_addr = R0_addr[25:0];
  assign mem_60_2_R0_clk = R0_clk;
  assign mem_60_2_R0_en = R0_en & R0_addr_sel == 8'h3c;
  assign mem_60_2_W0_addr = W0_addr[25:0];
  assign mem_60_2_W0_clk = W0_clk;
  assign mem_60_2_W0_data = W0_data[23:16];
  assign mem_60_2_W0_en = W0_en & W0_addr_sel == 8'h3c;
  assign mem_60_2_W0_mask = W0_mask[2];
  assign mem_60_3_R0_addr = R0_addr[25:0];
  assign mem_60_3_R0_clk = R0_clk;
  assign mem_60_3_R0_en = R0_en & R0_addr_sel == 8'h3c;
  assign mem_60_3_W0_addr = W0_addr[25:0];
  assign mem_60_3_W0_clk = W0_clk;
  assign mem_60_3_W0_data = W0_data[31:24];
  assign mem_60_3_W0_en = W0_en & W0_addr_sel == 8'h3c;
  assign mem_60_3_W0_mask = W0_mask[3];
  assign mem_60_4_R0_addr = R0_addr[25:0];
  assign mem_60_4_R0_clk = R0_clk;
  assign mem_60_4_R0_en = R0_en & R0_addr_sel == 8'h3c;
  assign mem_60_4_W0_addr = W0_addr[25:0];
  assign mem_60_4_W0_clk = W0_clk;
  assign mem_60_4_W0_data = W0_data[39:32];
  assign mem_60_4_W0_en = W0_en & W0_addr_sel == 8'h3c;
  assign mem_60_4_W0_mask = W0_mask[4];
  assign mem_60_5_R0_addr = R0_addr[25:0];
  assign mem_60_5_R0_clk = R0_clk;
  assign mem_60_5_R0_en = R0_en & R0_addr_sel == 8'h3c;
  assign mem_60_5_W0_addr = W0_addr[25:0];
  assign mem_60_5_W0_clk = W0_clk;
  assign mem_60_5_W0_data = W0_data[47:40];
  assign mem_60_5_W0_en = W0_en & W0_addr_sel == 8'h3c;
  assign mem_60_5_W0_mask = W0_mask[5];
  assign mem_60_6_R0_addr = R0_addr[25:0];
  assign mem_60_6_R0_clk = R0_clk;
  assign mem_60_6_R0_en = R0_en & R0_addr_sel == 8'h3c;
  assign mem_60_6_W0_addr = W0_addr[25:0];
  assign mem_60_6_W0_clk = W0_clk;
  assign mem_60_6_W0_data = W0_data[55:48];
  assign mem_60_6_W0_en = W0_en & W0_addr_sel == 8'h3c;
  assign mem_60_6_W0_mask = W0_mask[6];
  assign mem_60_7_R0_addr = R0_addr[25:0];
  assign mem_60_7_R0_clk = R0_clk;
  assign mem_60_7_R0_en = R0_en & R0_addr_sel == 8'h3c;
  assign mem_60_7_W0_addr = W0_addr[25:0];
  assign mem_60_7_W0_clk = W0_clk;
  assign mem_60_7_W0_data = W0_data[63:56];
  assign mem_60_7_W0_en = W0_en & W0_addr_sel == 8'h3c;
  assign mem_60_7_W0_mask = W0_mask[7];
  assign mem_61_0_R0_addr = R0_addr[25:0];
  assign mem_61_0_R0_clk = R0_clk;
  assign mem_61_0_R0_en = R0_en & R0_addr_sel == 8'h3d;
  assign mem_61_0_W0_addr = W0_addr[25:0];
  assign mem_61_0_W0_clk = W0_clk;
  assign mem_61_0_W0_data = W0_data[7:0];
  assign mem_61_0_W0_en = W0_en & W0_addr_sel == 8'h3d;
  assign mem_61_0_W0_mask = W0_mask[0];
  assign mem_61_1_R0_addr = R0_addr[25:0];
  assign mem_61_1_R0_clk = R0_clk;
  assign mem_61_1_R0_en = R0_en & R0_addr_sel == 8'h3d;
  assign mem_61_1_W0_addr = W0_addr[25:0];
  assign mem_61_1_W0_clk = W0_clk;
  assign mem_61_1_W0_data = W0_data[15:8];
  assign mem_61_1_W0_en = W0_en & W0_addr_sel == 8'h3d;
  assign mem_61_1_W0_mask = W0_mask[1];
  assign mem_61_2_R0_addr = R0_addr[25:0];
  assign mem_61_2_R0_clk = R0_clk;
  assign mem_61_2_R0_en = R0_en & R0_addr_sel == 8'h3d;
  assign mem_61_2_W0_addr = W0_addr[25:0];
  assign mem_61_2_W0_clk = W0_clk;
  assign mem_61_2_W0_data = W0_data[23:16];
  assign mem_61_2_W0_en = W0_en & W0_addr_sel == 8'h3d;
  assign mem_61_2_W0_mask = W0_mask[2];
  assign mem_61_3_R0_addr = R0_addr[25:0];
  assign mem_61_3_R0_clk = R0_clk;
  assign mem_61_3_R0_en = R0_en & R0_addr_sel == 8'h3d;
  assign mem_61_3_W0_addr = W0_addr[25:0];
  assign mem_61_3_W0_clk = W0_clk;
  assign mem_61_3_W0_data = W0_data[31:24];
  assign mem_61_3_W0_en = W0_en & W0_addr_sel == 8'h3d;
  assign mem_61_3_W0_mask = W0_mask[3];
  assign mem_61_4_R0_addr = R0_addr[25:0];
  assign mem_61_4_R0_clk = R0_clk;
  assign mem_61_4_R0_en = R0_en & R0_addr_sel == 8'h3d;
  assign mem_61_4_W0_addr = W0_addr[25:0];
  assign mem_61_4_W0_clk = W0_clk;
  assign mem_61_4_W0_data = W0_data[39:32];
  assign mem_61_4_W0_en = W0_en & W0_addr_sel == 8'h3d;
  assign mem_61_4_W0_mask = W0_mask[4];
  assign mem_61_5_R0_addr = R0_addr[25:0];
  assign mem_61_5_R0_clk = R0_clk;
  assign mem_61_5_R0_en = R0_en & R0_addr_sel == 8'h3d;
  assign mem_61_5_W0_addr = W0_addr[25:0];
  assign mem_61_5_W0_clk = W0_clk;
  assign mem_61_5_W0_data = W0_data[47:40];
  assign mem_61_5_W0_en = W0_en & W0_addr_sel == 8'h3d;
  assign mem_61_5_W0_mask = W0_mask[5];
  assign mem_61_6_R0_addr = R0_addr[25:0];
  assign mem_61_6_R0_clk = R0_clk;
  assign mem_61_6_R0_en = R0_en & R0_addr_sel == 8'h3d;
  assign mem_61_6_W0_addr = W0_addr[25:0];
  assign mem_61_6_W0_clk = W0_clk;
  assign mem_61_6_W0_data = W0_data[55:48];
  assign mem_61_6_W0_en = W0_en & W0_addr_sel == 8'h3d;
  assign mem_61_6_W0_mask = W0_mask[6];
  assign mem_61_7_R0_addr = R0_addr[25:0];
  assign mem_61_7_R0_clk = R0_clk;
  assign mem_61_7_R0_en = R0_en & R0_addr_sel == 8'h3d;
  assign mem_61_7_W0_addr = W0_addr[25:0];
  assign mem_61_7_W0_clk = W0_clk;
  assign mem_61_7_W0_data = W0_data[63:56];
  assign mem_61_7_W0_en = W0_en & W0_addr_sel == 8'h3d;
  assign mem_61_7_W0_mask = W0_mask[7];
  assign mem_62_0_R0_addr = R0_addr[25:0];
  assign mem_62_0_R0_clk = R0_clk;
  assign mem_62_0_R0_en = R0_en & R0_addr_sel == 8'h3e;
  assign mem_62_0_W0_addr = W0_addr[25:0];
  assign mem_62_0_W0_clk = W0_clk;
  assign mem_62_0_W0_data = W0_data[7:0];
  assign mem_62_0_W0_en = W0_en & W0_addr_sel == 8'h3e;
  assign mem_62_0_W0_mask = W0_mask[0];
  assign mem_62_1_R0_addr = R0_addr[25:0];
  assign mem_62_1_R0_clk = R0_clk;
  assign mem_62_1_R0_en = R0_en & R0_addr_sel == 8'h3e;
  assign mem_62_1_W0_addr = W0_addr[25:0];
  assign mem_62_1_W0_clk = W0_clk;
  assign mem_62_1_W0_data = W0_data[15:8];
  assign mem_62_1_W0_en = W0_en & W0_addr_sel == 8'h3e;
  assign mem_62_1_W0_mask = W0_mask[1];
  assign mem_62_2_R0_addr = R0_addr[25:0];
  assign mem_62_2_R0_clk = R0_clk;
  assign mem_62_2_R0_en = R0_en & R0_addr_sel == 8'h3e;
  assign mem_62_2_W0_addr = W0_addr[25:0];
  assign mem_62_2_W0_clk = W0_clk;
  assign mem_62_2_W0_data = W0_data[23:16];
  assign mem_62_2_W0_en = W0_en & W0_addr_sel == 8'h3e;
  assign mem_62_2_W0_mask = W0_mask[2];
  assign mem_62_3_R0_addr = R0_addr[25:0];
  assign mem_62_3_R0_clk = R0_clk;
  assign mem_62_3_R0_en = R0_en & R0_addr_sel == 8'h3e;
  assign mem_62_3_W0_addr = W0_addr[25:0];
  assign mem_62_3_W0_clk = W0_clk;
  assign mem_62_3_W0_data = W0_data[31:24];
  assign mem_62_3_W0_en = W0_en & W0_addr_sel == 8'h3e;
  assign mem_62_3_W0_mask = W0_mask[3];
  assign mem_62_4_R0_addr = R0_addr[25:0];
  assign mem_62_4_R0_clk = R0_clk;
  assign mem_62_4_R0_en = R0_en & R0_addr_sel == 8'h3e;
  assign mem_62_4_W0_addr = W0_addr[25:0];
  assign mem_62_4_W0_clk = W0_clk;
  assign mem_62_4_W0_data = W0_data[39:32];
  assign mem_62_4_W0_en = W0_en & W0_addr_sel == 8'h3e;
  assign mem_62_4_W0_mask = W0_mask[4];
  assign mem_62_5_R0_addr = R0_addr[25:0];
  assign mem_62_5_R0_clk = R0_clk;
  assign mem_62_5_R0_en = R0_en & R0_addr_sel == 8'h3e;
  assign mem_62_5_W0_addr = W0_addr[25:0];
  assign mem_62_5_W0_clk = W0_clk;
  assign mem_62_5_W0_data = W0_data[47:40];
  assign mem_62_5_W0_en = W0_en & W0_addr_sel == 8'h3e;
  assign mem_62_5_W0_mask = W0_mask[5];
  assign mem_62_6_R0_addr = R0_addr[25:0];
  assign mem_62_6_R0_clk = R0_clk;
  assign mem_62_6_R0_en = R0_en & R0_addr_sel == 8'h3e;
  assign mem_62_6_W0_addr = W0_addr[25:0];
  assign mem_62_6_W0_clk = W0_clk;
  assign mem_62_6_W0_data = W0_data[55:48];
  assign mem_62_6_W0_en = W0_en & W0_addr_sel == 8'h3e;
  assign mem_62_6_W0_mask = W0_mask[6];
  assign mem_62_7_R0_addr = R0_addr[25:0];
  assign mem_62_7_R0_clk = R0_clk;
  assign mem_62_7_R0_en = R0_en & R0_addr_sel == 8'h3e;
  assign mem_62_7_W0_addr = W0_addr[25:0];
  assign mem_62_7_W0_clk = W0_clk;
  assign mem_62_7_W0_data = W0_data[63:56];
  assign mem_62_7_W0_en = W0_en & W0_addr_sel == 8'h3e;
  assign mem_62_7_W0_mask = W0_mask[7];
  assign mem_63_0_R0_addr = R0_addr[25:0];
  assign mem_63_0_R0_clk = R0_clk;
  assign mem_63_0_R0_en = R0_en & R0_addr_sel == 8'h3f;
  assign mem_63_0_W0_addr = W0_addr[25:0];
  assign mem_63_0_W0_clk = W0_clk;
  assign mem_63_0_W0_data = W0_data[7:0];
  assign mem_63_0_W0_en = W0_en & W0_addr_sel == 8'h3f;
  assign mem_63_0_W0_mask = W0_mask[0];
  assign mem_63_1_R0_addr = R0_addr[25:0];
  assign mem_63_1_R0_clk = R0_clk;
  assign mem_63_1_R0_en = R0_en & R0_addr_sel == 8'h3f;
  assign mem_63_1_W0_addr = W0_addr[25:0];
  assign mem_63_1_W0_clk = W0_clk;
  assign mem_63_1_W0_data = W0_data[15:8];
  assign mem_63_1_W0_en = W0_en & W0_addr_sel == 8'h3f;
  assign mem_63_1_W0_mask = W0_mask[1];
  assign mem_63_2_R0_addr = R0_addr[25:0];
  assign mem_63_2_R0_clk = R0_clk;
  assign mem_63_2_R0_en = R0_en & R0_addr_sel == 8'h3f;
  assign mem_63_2_W0_addr = W0_addr[25:0];
  assign mem_63_2_W0_clk = W0_clk;
  assign mem_63_2_W0_data = W0_data[23:16];
  assign mem_63_2_W0_en = W0_en & W0_addr_sel == 8'h3f;
  assign mem_63_2_W0_mask = W0_mask[2];
  assign mem_63_3_R0_addr = R0_addr[25:0];
  assign mem_63_3_R0_clk = R0_clk;
  assign mem_63_3_R0_en = R0_en & R0_addr_sel == 8'h3f;
  assign mem_63_3_W0_addr = W0_addr[25:0];
  assign mem_63_3_W0_clk = W0_clk;
  assign mem_63_3_W0_data = W0_data[31:24];
  assign mem_63_3_W0_en = W0_en & W0_addr_sel == 8'h3f;
  assign mem_63_3_W0_mask = W0_mask[3];
  assign mem_63_4_R0_addr = R0_addr[25:0];
  assign mem_63_4_R0_clk = R0_clk;
  assign mem_63_4_R0_en = R0_en & R0_addr_sel == 8'h3f;
  assign mem_63_4_W0_addr = W0_addr[25:0];
  assign mem_63_4_W0_clk = W0_clk;
  assign mem_63_4_W0_data = W0_data[39:32];
  assign mem_63_4_W0_en = W0_en & W0_addr_sel == 8'h3f;
  assign mem_63_4_W0_mask = W0_mask[4];
  assign mem_63_5_R0_addr = R0_addr[25:0];
  assign mem_63_5_R0_clk = R0_clk;
  assign mem_63_5_R0_en = R0_en & R0_addr_sel == 8'h3f;
  assign mem_63_5_W0_addr = W0_addr[25:0];
  assign mem_63_5_W0_clk = W0_clk;
  assign mem_63_5_W0_data = W0_data[47:40];
  assign mem_63_5_W0_en = W0_en & W0_addr_sel == 8'h3f;
  assign mem_63_5_W0_mask = W0_mask[5];
  assign mem_63_6_R0_addr = R0_addr[25:0];
  assign mem_63_6_R0_clk = R0_clk;
  assign mem_63_6_R0_en = R0_en & R0_addr_sel == 8'h3f;
  assign mem_63_6_W0_addr = W0_addr[25:0];
  assign mem_63_6_W0_clk = W0_clk;
  assign mem_63_6_W0_data = W0_data[55:48];
  assign mem_63_6_W0_en = W0_en & W0_addr_sel == 8'h3f;
  assign mem_63_6_W0_mask = W0_mask[6];
  assign mem_63_7_R0_addr = R0_addr[25:0];
  assign mem_63_7_R0_clk = R0_clk;
  assign mem_63_7_R0_en = R0_en & R0_addr_sel == 8'h3f;
  assign mem_63_7_W0_addr = W0_addr[25:0];
  assign mem_63_7_W0_clk = W0_clk;
  assign mem_63_7_W0_data = W0_data[63:56];
  assign mem_63_7_W0_en = W0_en & W0_addr_sel == 8'h3f;
  assign mem_63_7_W0_mask = W0_mask[7];
  assign mem_64_0_R0_addr = R0_addr[25:0];
  assign mem_64_0_R0_clk = R0_clk;
  assign mem_64_0_R0_en = R0_en & R0_addr_sel == 8'h40;
  assign mem_64_0_W0_addr = W0_addr[25:0];
  assign mem_64_0_W0_clk = W0_clk;
  assign mem_64_0_W0_data = W0_data[7:0];
  assign mem_64_0_W0_en = W0_en & W0_addr_sel == 8'h40;
  assign mem_64_0_W0_mask = W0_mask[0];
  assign mem_64_1_R0_addr = R0_addr[25:0];
  assign mem_64_1_R0_clk = R0_clk;
  assign mem_64_1_R0_en = R0_en & R0_addr_sel == 8'h40;
  assign mem_64_1_W0_addr = W0_addr[25:0];
  assign mem_64_1_W0_clk = W0_clk;
  assign mem_64_1_W0_data = W0_data[15:8];
  assign mem_64_1_W0_en = W0_en & W0_addr_sel == 8'h40;
  assign mem_64_1_W0_mask = W0_mask[1];
  assign mem_64_2_R0_addr = R0_addr[25:0];
  assign mem_64_2_R0_clk = R0_clk;
  assign mem_64_2_R0_en = R0_en & R0_addr_sel == 8'h40;
  assign mem_64_2_W0_addr = W0_addr[25:0];
  assign mem_64_2_W0_clk = W0_clk;
  assign mem_64_2_W0_data = W0_data[23:16];
  assign mem_64_2_W0_en = W0_en & W0_addr_sel == 8'h40;
  assign mem_64_2_W0_mask = W0_mask[2];
  assign mem_64_3_R0_addr = R0_addr[25:0];
  assign mem_64_3_R0_clk = R0_clk;
  assign mem_64_3_R0_en = R0_en & R0_addr_sel == 8'h40;
  assign mem_64_3_W0_addr = W0_addr[25:0];
  assign mem_64_3_W0_clk = W0_clk;
  assign mem_64_3_W0_data = W0_data[31:24];
  assign mem_64_3_W0_en = W0_en & W0_addr_sel == 8'h40;
  assign mem_64_3_W0_mask = W0_mask[3];
  assign mem_64_4_R0_addr = R0_addr[25:0];
  assign mem_64_4_R0_clk = R0_clk;
  assign mem_64_4_R0_en = R0_en & R0_addr_sel == 8'h40;
  assign mem_64_4_W0_addr = W0_addr[25:0];
  assign mem_64_4_W0_clk = W0_clk;
  assign mem_64_4_W0_data = W0_data[39:32];
  assign mem_64_4_W0_en = W0_en & W0_addr_sel == 8'h40;
  assign mem_64_4_W0_mask = W0_mask[4];
  assign mem_64_5_R0_addr = R0_addr[25:0];
  assign mem_64_5_R0_clk = R0_clk;
  assign mem_64_5_R0_en = R0_en & R0_addr_sel == 8'h40;
  assign mem_64_5_W0_addr = W0_addr[25:0];
  assign mem_64_5_W0_clk = W0_clk;
  assign mem_64_5_W0_data = W0_data[47:40];
  assign mem_64_5_W0_en = W0_en & W0_addr_sel == 8'h40;
  assign mem_64_5_W0_mask = W0_mask[5];
  assign mem_64_6_R0_addr = R0_addr[25:0];
  assign mem_64_6_R0_clk = R0_clk;
  assign mem_64_6_R0_en = R0_en & R0_addr_sel == 8'h40;
  assign mem_64_6_W0_addr = W0_addr[25:0];
  assign mem_64_6_W0_clk = W0_clk;
  assign mem_64_6_W0_data = W0_data[55:48];
  assign mem_64_6_W0_en = W0_en & W0_addr_sel == 8'h40;
  assign mem_64_6_W0_mask = W0_mask[6];
  assign mem_64_7_R0_addr = R0_addr[25:0];
  assign mem_64_7_R0_clk = R0_clk;
  assign mem_64_7_R0_en = R0_en & R0_addr_sel == 8'h40;
  assign mem_64_7_W0_addr = W0_addr[25:0];
  assign mem_64_7_W0_clk = W0_clk;
  assign mem_64_7_W0_data = W0_data[63:56];
  assign mem_64_7_W0_en = W0_en & W0_addr_sel == 8'h40;
  assign mem_64_7_W0_mask = W0_mask[7];
  assign mem_65_0_R0_addr = R0_addr[25:0];
  assign mem_65_0_R0_clk = R0_clk;
  assign mem_65_0_R0_en = R0_en & R0_addr_sel == 8'h41;
  assign mem_65_0_W0_addr = W0_addr[25:0];
  assign mem_65_0_W0_clk = W0_clk;
  assign mem_65_0_W0_data = W0_data[7:0];
  assign mem_65_0_W0_en = W0_en & W0_addr_sel == 8'h41;
  assign mem_65_0_W0_mask = W0_mask[0];
  assign mem_65_1_R0_addr = R0_addr[25:0];
  assign mem_65_1_R0_clk = R0_clk;
  assign mem_65_1_R0_en = R0_en & R0_addr_sel == 8'h41;
  assign mem_65_1_W0_addr = W0_addr[25:0];
  assign mem_65_1_W0_clk = W0_clk;
  assign mem_65_1_W0_data = W0_data[15:8];
  assign mem_65_1_W0_en = W0_en & W0_addr_sel == 8'h41;
  assign mem_65_1_W0_mask = W0_mask[1];
  assign mem_65_2_R0_addr = R0_addr[25:0];
  assign mem_65_2_R0_clk = R0_clk;
  assign mem_65_2_R0_en = R0_en & R0_addr_sel == 8'h41;
  assign mem_65_2_W0_addr = W0_addr[25:0];
  assign mem_65_2_W0_clk = W0_clk;
  assign mem_65_2_W0_data = W0_data[23:16];
  assign mem_65_2_W0_en = W0_en & W0_addr_sel == 8'h41;
  assign mem_65_2_W0_mask = W0_mask[2];
  assign mem_65_3_R0_addr = R0_addr[25:0];
  assign mem_65_3_R0_clk = R0_clk;
  assign mem_65_3_R0_en = R0_en & R0_addr_sel == 8'h41;
  assign mem_65_3_W0_addr = W0_addr[25:0];
  assign mem_65_3_W0_clk = W0_clk;
  assign mem_65_3_W0_data = W0_data[31:24];
  assign mem_65_3_W0_en = W0_en & W0_addr_sel == 8'h41;
  assign mem_65_3_W0_mask = W0_mask[3];
  assign mem_65_4_R0_addr = R0_addr[25:0];
  assign mem_65_4_R0_clk = R0_clk;
  assign mem_65_4_R0_en = R0_en & R0_addr_sel == 8'h41;
  assign mem_65_4_W0_addr = W0_addr[25:0];
  assign mem_65_4_W0_clk = W0_clk;
  assign mem_65_4_W0_data = W0_data[39:32];
  assign mem_65_4_W0_en = W0_en & W0_addr_sel == 8'h41;
  assign mem_65_4_W0_mask = W0_mask[4];
  assign mem_65_5_R0_addr = R0_addr[25:0];
  assign mem_65_5_R0_clk = R0_clk;
  assign mem_65_5_R0_en = R0_en & R0_addr_sel == 8'h41;
  assign mem_65_5_W0_addr = W0_addr[25:0];
  assign mem_65_5_W0_clk = W0_clk;
  assign mem_65_5_W0_data = W0_data[47:40];
  assign mem_65_5_W0_en = W0_en & W0_addr_sel == 8'h41;
  assign mem_65_5_W0_mask = W0_mask[5];
  assign mem_65_6_R0_addr = R0_addr[25:0];
  assign mem_65_6_R0_clk = R0_clk;
  assign mem_65_6_R0_en = R0_en & R0_addr_sel == 8'h41;
  assign mem_65_6_W0_addr = W0_addr[25:0];
  assign mem_65_6_W0_clk = W0_clk;
  assign mem_65_6_W0_data = W0_data[55:48];
  assign mem_65_6_W0_en = W0_en & W0_addr_sel == 8'h41;
  assign mem_65_6_W0_mask = W0_mask[6];
  assign mem_65_7_R0_addr = R0_addr[25:0];
  assign mem_65_7_R0_clk = R0_clk;
  assign mem_65_7_R0_en = R0_en & R0_addr_sel == 8'h41;
  assign mem_65_7_W0_addr = W0_addr[25:0];
  assign mem_65_7_W0_clk = W0_clk;
  assign mem_65_7_W0_data = W0_data[63:56];
  assign mem_65_7_W0_en = W0_en & W0_addr_sel == 8'h41;
  assign mem_65_7_W0_mask = W0_mask[7];
  assign mem_66_0_R0_addr = R0_addr[25:0];
  assign mem_66_0_R0_clk = R0_clk;
  assign mem_66_0_R0_en = R0_en & R0_addr_sel == 8'h42;
  assign mem_66_0_W0_addr = W0_addr[25:0];
  assign mem_66_0_W0_clk = W0_clk;
  assign mem_66_0_W0_data = W0_data[7:0];
  assign mem_66_0_W0_en = W0_en & W0_addr_sel == 8'h42;
  assign mem_66_0_W0_mask = W0_mask[0];
  assign mem_66_1_R0_addr = R0_addr[25:0];
  assign mem_66_1_R0_clk = R0_clk;
  assign mem_66_1_R0_en = R0_en & R0_addr_sel == 8'h42;
  assign mem_66_1_W0_addr = W0_addr[25:0];
  assign mem_66_1_W0_clk = W0_clk;
  assign mem_66_1_W0_data = W0_data[15:8];
  assign mem_66_1_W0_en = W0_en & W0_addr_sel == 8'h42;
  assign mem_66_1_W0_mask = W0_mask[1];
  assign mem_66_2_R0_addr = R0_addr[25:0];
  assign mem_66_2_R0_clk = R0_clk;
  assign mem_66_2_R0_en = R0_en & R0_addr_sel == 8'h42;
  assign mem_66_2_W0_addr = W0_addr[25:0];
  assign mem_66_2_W0_clk = W0_clk;
  assign mem_66_2_W0_data = W0_data[23:16];
  assign mem_66_2_W0_en = W0_en & W0_addr_sel == 8'h42;
  assign mem_66_2_W0_mask = W0_mask[2];
  assign mem_66_3_R0_addr = R0_addr[25:0];
  assign mem_66_3_R0_clk = R0_clk;
  assign mem_66_3_R0_en = R0_en & R0_addr_sel == 8'h42;
  assign mem_66_3_W0_addr = W0_addr[25:0];
  assign mem_66_3_W0_clk = W0_clk;
  assign mem_66_3_W0_data = W0_data[31:24];
  assign mem_66_3_W0_en = W0_en & W0_addr_sel == 8'h42;
  assign mem_66_3_W0_mask = W0_mask[3];
  assign mem_66_4_R0_addr = R0_addr[25:0];
  assign mem_66_4_R0_clk = R0_clk;
  assign mem_66_4_R0_en = R0_en & R0_addr_sel == 8'h42;
  assign mem_66_4_W0_addr = W0_addr[25:0];
  assign mem_66_4_W0_clk = W0_clk;
  assign mem_66_4_W0_data = W0_data[39:32];
  assign mem_66_4_W0_en = W0_en & W0_addr_sel == 8'h42;
  assign mem_66_4_W0_mask = W0_mask[4];
  assign mem_66_5_R0_addr = R0_addr[25:0];
  assign mem_66_5_R0_clk = R0_clk;
  assign mem_66_5_R0_en = R0_en & R0_addr_sel == 8'h42;
  assign mem_66_5_W0_addr = W0_addr[25:0];
  assign mem_66_5_W0_clk = W0_clk;
  assign mem_66_5_W0_data = W0_data[47:40];
  assign mem_66_5_W0_en = W0_en & W0_addr_sel == 8'h42;
  assign mem_66_5_W0_mask = W0_mask[5];
  assign mem_66_6_R0_addr = R0_addr[25:0];
  assign mem_66_6_R0_clk = R0_clk;
  assign mem_66_6_R0_en = R0_en & R0_addr_sel == 8'h42;
  assign mem_66_6_W0_addr = W0_addr[25:0];
  assign mem_66_6_W0_clk = W0_clk;
  assign mem_66_6_W0_data = W0_data[55:48];
  assign mem_66_6_W0_en = W0_en & W0_addr_sel == 8'h42;
  assign mem_66_6_W0_mask = W0_mask[6];
  assign mem_66_7_R0_addr = R0_addr[25:0];
  assign mem_66_7_R0_clk = R0_clk;
  assign mem_66_7_R0_en = R0_en & R0_addr_sel == 8'h42;
  assign mem_66_7_W0_addr = W0_addr[25:0];
  assign mem_66_7_W0_clk = W0_clk;
  assign mem_66_7_W0_data = W0_data[63:56];
  assign mem_66_7_W0_en = W0_en & W0_addr_sel == 8'h42;
  assign mem_66_7_W0_mask = W0_mask[7];
  assign mem_67_0_R0_addr = R0_addr[25:0];
  assign mem_67_0_R0_clk = R0_clk;
  assign mem_67_0_R0_en = R0_en & R0_addr_sel == 8'h43;
  assign mem_67_0_W0_addr = W0_addr[25:0];
  assign mem_67_0_W0_clk = W0_clk;
  assign mem_67_0_W0_data = W0_data[7:0];
  assign mem_67_0_W0_en = W0_en & W0_addr_sel == 8'h43;
  assign mem_67_0_W0_mask = W0_mask[0];
  assign mem_67_1_R0_addr = R0_addr[25:0];
  assign mem_67_1_R0_clk = R0_clk;
  assign mem_67_1_R0_en = R0_en & R0_addr_sel == 8'h43;
  assign mem_67_1_W0_addr = W0_addr[25:0];
  assign mem_67_1_W0_clk = W0_clk;
  assign mem_67_1_W0_data = W0_data[15:8];
  assign mem_67_1_W0_en = W0_en & W0_addr_sel == 8'h43;
  assign mem_67_1_W0_mask = W0_mask[1];
  assign mem_67_2_R0_addr = R0_addr[25:0];
  assign mem_67_2_R0_clk = R0_clk;
  assign mem_67_2_R0_en = R0_en & R0_addr_sel == 8'h43;
  assign mem_67_2_W0_addr = W0_addr[25:0];
  assign mem_67_2_W0_clk = W0_clk;
  assign mem_67_2_W0_data = W0_data[23:16];
  assign mem_67_2_W0_en = W0_en & W0_addr_sel == 8'h43;
  assign mem_67_2_W0_mask = W0_mask[2];
  assign mem_67_3_R0_addr = R0_addr[25:0];
  assign mem_67_3_R0_clk = R0_clk;
  assign mem_67_3_R0_en = R0_en & R0_addr_sel == 8'h43;
  assign mem_67_3_W0_addr = W0_addr[25:0];
  assign mem_67_3_W0_clk = W0_clk;
  assign mem_67_3_W0_data = W0_data[31:24];
  assign mem_67_3_W0_en = W0_en & W0_addr_sel == 8'h43;
  assign mem_67_3_W0_mask = W0_mask[3];
  assign mem_67_4_R0_addr = R0_addr[25:0];
  assign mem_67_4_R0_clk = R0_clk;
  assign mem_67_4_R0_en = R0_en & R0_addr_sel == 8'h43;
  assign mem_67_4_W0_addr = W0_addr[25:0];
  assign mem_67_4_W0_clk = W0_clk;
  assign mem_67_4_W0_data = W0_data[39:32];
  assign mem_67_4_W0_en = W0_en & W0_addr_sel == 8'h43;
  assign mem_67_4_W0_mask = W0_mask[4];
  assign mem_67_5_R0_addr = R0_addr[25:0];
  assign mem_67_5_R0_clk = R0_clk;
  assign mem_67_5_R0_en = R0_en & R0_addr_sel == 8'h43;
  assign mem_67_5_W0_addr = W0_addr[25:0];
  assign mem_67_5_W0_clk = W0_clk;
  assign mem_67_5_W0_data = W0_data[47:40];
  assign mem_67_5_W0_en = W0_en & W0_addr_sel == 8'h43;
  assign mem_67_5_W0_mask = W0_mask[5];
  assign mem_67_6_R0_addr = R0_addr[25:0];
  assign mem_67_6_R0_clk = R0_clk;
  assign mem_67_6_R0_en = R0_en & R0_addr_sel == 8'h43;
  assign mem_67_6_W0_addr = W0_addr[25:0];
  assign mem_67_6_W0_clk = W0_clk;
  assign mem_67_6_W0_data = W0_data[55:48];
  assign mem_67_6_W0_en = W0_en & W0_addr_sel == 8'h43;
  assign mem_67_6_W0_mask = W0_mask[6];
  assign mem_67_7_R0_addr = R0_addr[25:0];
  assign mem_67_7_R0_clk = R0_clk;
  assign mem_67_7_R0_en = R0_en & R0_addr_sel == 8'h43;
  assign mem_67_7_W0_addr = W0_addr[25:0];
  assign mem_67_7_W0_clk = W0_clk;
  assign mem_67_7_W0_data = W0_data[63:56];
  assign mem_67_7_W0_en = W0_en & W0_addr_sel == 8'h43;
  assign mem_67_7_W0_mask = W0_mask[7];
  assign mem_68_0_R0_addr = R0_addr[25:0];
  assign mem_68_0_R0_clk = R0_clk;
  assign mem_68_0_R0_en = R0_en & R0_addr_sel == 8'h44;
  assign mem_68_0_W0_addr = W0_addr[25:0];
  assign mem_68_0_W0_clk = W0_clk;
  assign mem_68_0_W0_data = W0_data[7:0];
  assign mem_68_0_W0_en = W0_en & W0_addr_sel == 8'h44;
  assign mem_68_0_W0_mask = W0_mask[0];
  assign mem_68_1_R0_addr = R0_addr[25:0];
  assign mem_68_1_R0_clk = R0_clk;
  assign mem_68_1_R0_en = R0_en & R0_addr_sel == 8'h44;
  assign mem_68_1_W0_addr = W0_addr[25:0];
  assign mem_68_1_W0_clk = W0_clk;
  assign mem_68_1_W0_data = W0_data[15:8];
  assign mem_68_1_W0_en = W0_en & W0_addr_sel == 8'h44;
  assign mem_68_1_W0_mask = W0_mask[1];
  assign mem_68_2_R0_addr = R0_addr[25:0];
  assign mem_68_2_R0_clk = R0_clk;
  assign mem_68_2_R0_en = R0_en & R0_addr_sel == 8'h44;
  assign mem_68_2_W0_addr = W0_addr[25:0];
  assign mem_68_2_W0_clk = W0_clk;
  assign mem_68_2_W0_data = W0_data[23:16];
  assign mem_68_2_W0_en = W0_en & W0_addr_sel == 8'h44;
  assign mem_68_2_W0_mask = W0_mask[2];
  assign mem_68_3_R0_addr = R0_addr[25:0];
  assign mem_68_3_R0_clk = R0_clk;
  assign mem_68_3_R0_en = R0_en & R0_addr_sel == 8'h44;
  assign mem_68_3_W0_addr = W0_addr[25:0];
  assign mem_68_3_W0_clk = W0_clk;
  assign mem_68_3_W0_data = W0_data[31:24];
  assign mem_68_3_W0_en = W0_en & W0_addr_sel == 8'h44;
  assign mem_68_3_W0_mask = W0_mask[3];
  assign mem_68_4_R0_addr = R0_addr[25:0];
  assign mem_68_4_R0_clk = R0_clk;
  assign mem_68_4_R0_en = R0_en & R0_addr_sel == 8'h44;
  assign mem_68_4_W0_addr = W0_addr[25:0];
  assign mem_68_4_W0_clk = W0_clk;
  assign mem_68_4_W0_data = W0_data[39:32];
  assign mem_68_4_W0_en = W0_en & W0_addr_sel == 8'h44;
  assign mem_68_4_W0_mask = W0_mask[4];
  assign mem_68_5_R0_addr = R0_addr[25:0];
  assign mem_68_5_R0_clk = R0_clk;
  assign mem_68_5_R0_en = R0_en & R0_addr_sel == 8'h44;
  assign mem_68_5_W0_addr = W0_addr[25:0];
  assign mem_68_5_W0_clk = W0_clk;
  assign mem_68_5_W0_data = W0_data[47:40];
  assign mem_68_5_W0_en = W0_en & W0_addr_sel == 8'h44;
  assign mem_68_5_W0_mask = W0_mask[5];
  assign mem_68_6_R0_addr = R0_addr[25:0];
  assign mem_68_6_R0_clk = R0_clk;
  assign mem_68_6_R0_en = R0_en & R0_addr_sel == 8'h44;
  assign mem_68_6_W0_addr = W0_addr[25:0];
  assign mem_68_6_W0_clk = W0_clk;
  assign mem_68_6_W0_data = W0_data[55:48];
  assign mem_68_6_W0_en = W0_en & W0_addr_sel == 8'h44;
  assign mem_68_6_W0_mask = W0_mask[6];
  assign mem_68_7_R0_addr = R0_addr[25:0];
  assign mem_68_7_R0_clk = R0_clk;
  assign mem_68_7_R0_en = R0_en & R0_addr_sel == 8'h44;
  assign mem_68_7_W0_addr = W0_addr[25:0];
  assign mem_68_7_W0_clk = W0_clk;
  assign mem_68_7_W0_data = W0_data[63:56];
  assign mem_68_7_W0_en = W0_en & W0_addr_sel == 8'h44;
  assign mem_68_7_W0_mask = W0_mask[7];
  assign mem_69_0_R0_addr = R0_addr[25:0];
  assign mem_69_0_R0_clk = R0_clk;
  assign mem_69_0_R0_en = R0_en & R0_addr_sel == 8'h45;
  assign mem_69_0_W0_addr = W0_addr[25:0];
  assign mem_69_0_W0_clk = W0_clk;
  assign mem_69_0_W0_data = W0_data[7:0];
  assign mem_69_0_W0_en = W0_en & W0_addr_sel == 8'h45;
  assign mem_69_0_W0_mask = W0_mask[0];
  assign mem_69_1_R0_addr = R0_addr[25:0];
  assign mem_69_1_R0_clk = R0_clk;
  assign mem_69_1_R0_en = R0_en & R0_addr_sel == 8'h45;
  assign mem_69_1_W0_addr = W0_addr[25:0];
  assign mem_69_1_W0_clk = W0_clk;
  assign mem_69_1_W0_data = W0_data[15:8];
  assign mem_69_1_W0_en = W0_en & W0_addr_sel == 8'h45;
  assign mem_69_1_W0_mask = W0_mask[1];
  assign mem_69_2_R0_addr = R0_addr[25:0];
  assign mem_69_2_R0_clk = R0_clk;
  assign mem_69_2_R0_en = R0_en & R0_addr_sel == 8'h45;
  assign mem_69_2_W0_addr = W0_addr[25:0];
  assign mem_69_2_W0_clk = W0_clk;
  assign mem_69_2_W0_data = W0_data[23:16];
  assign mem_69_2_W0_en = W0_en & W0_addr_sel == 8'h45;
  assign mem_69_2_W0_mask = W0_mask[2];
  assign mem_69_3_R0_addr = R0_addr[25:0];
  assign mem_69_3_R0_clk = R0_clk;
  assign mem_69_3_R0_en = R0_en & R0_addr_sel == 8'h45;
  assign mem_69_3_W0_addr = W0_addr[25:0];
  assign mem_69_3_W0_clk = W0_clk;
  assign mem_69_3_W0_data = W0_data[31:24];
  assign mem_69_3_W0_en = W0_en & W0_addr_sel == 8'h45;
  assign mem_69_3_W0_mask = W0_mask[3];
  assign mem_69_4_R0_addr = R0_addr[25:0];
  assign mem_69_4_R0_clk = R0_clk;
  assign mem_69_4_R0_en = R0_en & R0_addr_sel == 8'h45;
  assign mem_69_4_W0_addr = W0_addr[25:0];
  assign mem_69_4_W0_clk = W0_clk;
  assign mem_69_4_W0_data = W0_data[39:32];
  assign mem_69_4_W0_en = W0_en & W0_addr_sel == 8'h45;
  assign mem_69_4_W0_mask = W0_mask[4];
  assign mem_69_5_R0_addr = R0_addr[25:0];
  assign mem_69_5_R0_clk = R0_clk;
  assign mem_69_5_R0_en = R0_en & R0_addr_sel == 8'h45;
  assign mem_69_5_W0_addr = W0_addr[25:0];
  assign mem_69_5_W0_clk = W0_clk;
  assign mem_69_5_W0_data = W0_data[47:40];
  assign mem_69_5_W0_en = W0_en & W0_addr_sel == 8'h45;
  assign mem_69_5_W0_mask = W0_mask[5];
  assign mem_69_6_R0_addr = R0_addr[25:0];
  assign mem_69_6_R0_clk = R0_clk;
  assign mem_69_6_R0_en = R0_en & R0_addr_sel == 8'h45;
  assign mem_69_6_W0_addr = W0_addr[25:0];
  assign mem_69_6_W0_clk = W0_clk;
  assign mem_69_6_W0_data = W0_data[55:48];
  assign mem_69_6_W0_en = W0_en & W0_addr_sel == 8'h45;
  assign mem_69_6_W0_mask = W0_mask[6];
  assign mem_69_7_R0_addr = R0_addr[25:0];
  assign mem_69_7_R0_clk = R0_clk;
  assign mem_69_7_R0_en = R0_en & R0_addr_sel == 8'h45;
  assign mem_69_7_W0_addr = W0_addr[25:0];
  assign mem_69_7_W0_clk = W0_clk;
  assign mem_69_7_W0_data = W0_data[63:56];
  assign mem_69_7_W0_en = W0_en & W0_addr_sel == 8'h45;
  assign mem_69_7_W0_mask = W0_mask[7];
  assign mem_70_0_R0_addr = R0_addr[25:0];
  assign mem_70_0_R0_clk = R0_clk;
  assign mem_70_0_R0_en = R0_en & R0_addr_sel == 8'h46;
  assign mem_70_0_W0_addr = W0_addr[25:0];
  assign mem_70_0_W0_clk = W0_clk;
  assign mem_70_0_W0_data = W0_data[7:0];
  assign mem_70_0_W0_en = W0_en & W0_addr_sel == 8'h46;
  assign mem_70_0_W0_mask = W0_mask[0];
  assign mem_70_1_R0_addr = R0_addr[25:0];
  assign mem_70_1_R0_clk = R0_clk;
  assign mem_70_1_R0_en = R0_en & R0_addr_sel == 8'h46;
  assign mem_70_1_W0_addr = W0_addr[25:0];
  assign mem_70_1_W0_clk = W0_clk;
  assign mem_70_1_W0_data = W0_data[15:8];
  assign mem_70_1_W0_en = W0_en & W0_addr_sel == 8'h46;
  assign mem_70_1_W0_mask = W0_mask[1];
  assign mem_70_2_R0_addr = R0_addr[25:0];
  assign mem_70_2_R0_clk = R0_clk;
  assign mem_70_2_R0_en = R0_en & R0_addr_sel == 8'h46;
  assign mem_70_2_W0_addr = W0_addr[25:0];
  assign mem_70_2_W0_clk = W0_clk;
  assign mem_70_2_W0_data = W0_data[23:16];
  assign mem_70_2_W0_en = W0_en & W0_addr_sel == 8'h46;
  assign mem_70_2_W0_mask = W0_mask[2];
  assign mem_70_3_R0_addr = R0_addr[25:0];
  assign mem_70_3_R0_clk = R0_clk;
  assign mem_70_3_R0_en = R0_en & R0_addr_sel == 8'h46;
  assign mem_70_3_W0_addr = W0_addr[25:0];
  assign mem_70_3_W0_clk = W0_clk;
  assign mem_70_3_W0_data = W0_data[31:24];
  assign mem_70_3_W0_en = W0_en & W0_addr_sel == 8'h46;
  assign mem_70_3_W0_mask = W0_mask[3];
  assign mem_70_4_R0_addr = R0_addr[25:0];
  assign mem_70_4_R0_clk = R0_clk;
  assign mem_70_4_R0_en = R0_en & R0_addr_sel == 8'h46;
  assign mem_70_4_W0_addr = W0_addr[25:0];
  assign mem_70_4_W0_clk = W0_clk;
  assign mem_70_4_W0_data = W0_data[39:32];
  assign mem_70_4_W0_en = W0_en & W0_addr_sel == 8'h46;
  assign mem_70_4_W0_mask = W0_mask[4];
  assign mem_70_5_R0_addr = R0_addr[25:0];
  assign mem_70_5_R0_clk = R0_clk;
  assign mem_70_5_R0_en = R0_en & R0_addr_sel == 8'h46;
  assign mem_70_5_W0_addr = W0_addr[25:0];
  assign mem_70_5_W0_clk = W0_clk;
  assign mem_70_5_W0_data = W0_data[47:40];
  assign mem_70_5_W0_en = W0_en & W0_addr_sel == 8'h46;
  assign mem_70_5_W0_mask = W0_mask[5];
  assign mem_70_6_R0_addr = R0_addr[25:0];
  assign mem_70_6_R0_clk = R0_clk;
  assign mem_70_6_R0_en = R0_en & R0_addr_sel == 8'h46;
  assign mem_70_6_W0_addr = W0_addr[25:0];
  assign mem_70_6_W0_clk = W0_clk;
  assign mem_70_6_W0_data = W0_data[55:48];
  assign mem_70_6_W0_en = W0_en & W0_addr_sel == 8'h46;
  assign mem_70_6_W0_mask = W0_mask[6];
  assign mem_70_7_R0_addr = R0_addr[25:0];
  assign mem_70_7_R0_clk = R0_clk;
  assign mem_70_7_R0_en = R0_en & R0_addr_sel == 8'h46;
  assign mem_70_7_W0_addr = W0_addr[25:0];
  assign mem_70_7_W0_clk = W0_clk;
  assign mem_70_7_W0_data = W0_data[63:56];
  assign mem_70_7_W0_en = W0_en & W0_addr_sel == 8'h46;
  assign mem_70_7_W0_mask = W0_mask[7];
  assign mem_71_0_R0_addr = R0_addr[25:0];
  assign mem_71_0_R0_clk = R0_clk;
  assign mem_71_0_R0_en = R0_en & R0_addr_sel == 8'h47;
  assign mem_71_0_W0_addr = W0_addr[25:0];
  assign mem_71_0_W0_clk = W0_clk;
  assign mem_71_0_W0_data = W0_data[7:0];
  assign mem_71_0_W0_en = W0_en & W0_addr_sel == 8'h47;
  assign mem_71_0_W0_mask = W0_mask[0];
  assign mem_71_1_R0_addr = R0_addr[25:0];
  assign mem_71_1_R0_clk = R0_clk;
  assign mem_71_1_R0_en = R0_en & R0_addr_sel == 8'h47;
  assign mem_71_1_W0_addr = W0_addr[25:0];
  assign mem_71_1_W0_clk = W0_clk;
  assign mem_71_1_W0_data = W0_data[15:8];
  assign mem_71_1_W0_en = W0_en & W0_addr_sel == 8'h47;
  assign mem_71_1_W0_mask = W0_mask[1];
  assign mem_71_2_R0_addr = R0_addr[25:0];
  assign mem_71_2_R0_clk = R0_clk;
  assign mem_71_2_R0_en = R0_en & R0_addr_sel == 8'h47;
  assign mem_71_2_W0_addr = W0_addr[25:0];
  assign mem_71_2_W0_clk = W0_clk;
  assign mem_71_2_W0_data = W0_data[23:16];
  assign mem_71_2_W0_en = W0_en & W0_addr_sel == 8'h47;
  assign mem_71_2_W0_mask = W0_mask[2];
  assign mem_71_3_R0_addr = R0_addr[25:0];
  assign mem_71_3_R0_clk = R0_clk;
  assign mem_71_3_R0_en = R0_en & R0_addr_sel == 8'h47;
  assign mem_71_3_W0_addr = W0_addr[25:0];
  assign mem_71_3_W0_clk = W0_clk;
  assign mem_71_3_W0_data = W0_data[31:24];
  assign mem_71_3_W0_en = W0_en & W0_addr_sel == 8'h47;
  assign mem_71_3_W0_mask = W0_mask[3];
  assign mem_71_4_R0_addr = R0_addr[25:0];
  assign mem_71_4_R0_clk = R0_clk;
  assign mem_71_4_R0_en = R0_en & R0_addr_sel == 8'h47;
  assign mem_71_4_W0_addr = W0_addr[25:0];
  assign mem_71_4_W0_clk = W0_clk;
  assign mem_71_4_W0_data = W0_data[39:32];
  assign mem_71_4_W0_en = W0_en & W0_addr_sel == 8'h47;
  assign mem_71_4_W0_mask = W0_mask[4];
  assign mem_71_5_R0_addr = R0_addr[25:0];
  assign mem_71_5_R0_clk = R0_clk;
  assign mem_71_5_R0_en = R0_en & R0_addr_sel == 8'h47;
  assign mem_71_5_W0_addr = W0_addr[25:0];
  assign mem_71_5_W0_clk = W0_clk;
  assign mem_71_5_W0_data = W0_data[47:40];
  assign mem_71_5_W0_en = W0_en & W0_addr_sel == 8'h47;
  assign mem_71_5_W0_mask = W0_mask[5];
  assign mem_71_6_R0_addr = R0_addr[25:0];
  assign mem_71_6_R0_clk = R0_clk;
  assign mem_71_6_R0_en = R0_en & R0_addr_sel == 8'h47;
  assign mem_71_6_W0_addr = W0_addr[25:0];
  assign mem_71_6_W0_clk = W0_clk;
  assign mem_71_6_W0_data = W0_data[55:48];
  assign mem_71_6_W0_en = W0_en & W0_addr_sel == 8'h47;
  assign mem_71_6_W0_mask = W0_mask[6];
  assign mem_71_7_R0_addr = R0_addr[25:0];
  assign mem_71_7_R0_clk = R0_clk;
  assign mem_71_7_R0_en = R0_en & R0_addr_sel == 8'h47;
  assign mem_71_7_W0_addr = W0_addr[25:0];
  assign mem_71_7_W0_clk = W0_clk;
  assign mem_71_7_W0_data = W0_data[63:56];
  assign mem_71_7_W0_en = W0_en & W0_addr_sel == 8'h47;
  assign mem_71_7_W0_mask = W0_mask[7];
  assign mem_72_0_R0_addr = R0_addr[25:0];
  assign mem_72_0_R0_clk = R0_clk;
  assign mem_72_0_R0_en = R0_en & R0_addr_sel == 8'h48;
  assign mem_72_0_W0_addr = W0_addr[25:0];
  assign mem_72_0_W0_clk = W0_clk;
  assign mem_72_0_W0_data = W0_data[7:0];
  assign mem_72_0_W0_en = W0_en & W0_addr_sel == 8'h48;
  assign mem_72_0_W0_mask = W0_mask[0];
  assign mem_72_1_R0_addr = R0_addr[25:0];
  assign mem_72_1_R0_clk = R0_clk;
  assign mem_72_1_R0_en = R0_en & R0_addr_sel == 8'h48;
  assign mem_72_1_W0_addr = W0_addr[25:0];
  assign mem_72_1_W0_clk = W0_clk;
  assign mem_72_1_W0_data = W0_data[15:8];
  assign mem_72_1_W0_en = W0_en & W0_addr_sel == 8'h48;
  assign mem_72_1_W0_mask = W0_mask[1];
  assign mem_72_2_R0_addr = R0_addr[25:0];
  assign mem_72_2_R0_clk = R0_clk;
  assign mem_72_2_R0_en = R0_en & R0_addr_sel == 8'h48;
  assign mem_72_2_W0_addr = W0_addr[25:0];
  assign mem_72_2_W0_clk = W0_clk;
  assign mem_72_2_W0_data = W0_data[23:16];
  assign mem_72_2_W0_en = W0_en & W0_addr_sel == 8'h48;
  assign mem_72_2_W0_mask = W0_mask[2];
  assign mem_72_3_R0_addr = R0_addr[25:0];
  assign mem_72_3_R0_clk = R0_clk;
  assign mem_72_3_R0_en = R0_en & R0_addr_sel == 8'h48;
  assign mem_72_3_W0_addr = W0_addr[25:0];
  assign mem_72_3_W0_clk = W0_clk;
  assign mem_72_3_W0_data = W0_data[31:24];
  assign mem_72_3_W0_en = W0_en & W0_addr_sel == 8'h48;
  assign mem_72_3_W0_mask = W0_mask[3];
  assign mem_72_4_R0_addr = R0_addr[25:0];
  assign mem_72_4_R0_clk = R0_clk;
  assign mem_72_4_R0_en = R0_en & R0_addr_sel == 8'h48;
  assign mem_72_4_W0_addr = W0_addr[25:0];
  assign mem_72_4_W0_clk = W0_clk;
  assign mem_72_4_W0_data = W0_data[39:32];
  assign mem_72_4_W0_en = W0_en & W0_addr_sel == 8'h48;
  assign mem_72_4_W0_mask = W0_mask[4];
  assign mem_72_5_R0_addr = R0_addr[25:0];
  assign mem_72_5_R0_clk = R0_clk;
  assign mem_72_5_R0_en = R0_en & R0_addr_sel == 8'h48;
  assign mem_72_5_W0_addr = W0_addr[25:0];
  assign mem_72_5_W0_clk = W0_clk;
  assign mem_72_5_W0_data = W0_data[47:40];
  assign mem_72_5_W0_en = W0_en & W0_addr_sel == 8'h48;
  assign mem_72_5_W0_mask = W0_mask[5];
  assign mem_72_6_R0_addr = R0_addr[25:0];
  assign mem_72_6_R0_clk = R0_clk;
  assign mem_72_6_R0_en = R0_en & R0_addr_sel == 8'h48;
  assign mem_72_6_W0_addr = W0_addr[25:0];
  assign mem_72_6_W0_clk = W0_clk;
  assign mem_72_6_W0_data = W0_data[55:48];
  assign mem_72_6_W0_en = W0_en & W0_addr_sel == 8'h48;
  assign mem_72_6_W0_mask = W0_mask[6];
  assign mem_72_7_R0_addr = R0_addr[25:0];
  assign mem_72_7_R0_clk = R0_clk;
  assign mem_72_7_R0_en = R0_en & R0_addr_sel == 8'h48;
  assign mem_72_7_W0_addr = W0_addr[25:0];
  assign mem_72_7_W0_clk = W0_clk;
  assign mem_72_7_W0_data = W0_data[63:56];
  assign mem_72_7_W0_en = W0_en & W0_addr_sel == 8'h48;
  assign mem_72_7_W0_mask = W0_mask[7];
  assign mem_73_0_R0_addr = R0_addr[25:0];
  assign mem_73_0_R0_clk = R0_clk;
  assign mem_73_0_R0_en = R0_en & R0_addr_sel == 8'h49;
  assign mem_73_0_W0_addr = W0_addr[25:0];
  assign mem_73_0_W0_clk = W0_clk;
  assign mem_73_0_W0_data = W0_data[7:0];
  assign mem_73_0_W0_en = W0_en & W0_addr_sel == 8'h49;
  assign mem_73_0_W0_mask = W0_mask[0];
  assign mem_73_1_R0_addr = R0_addr[25:0];
  assign mem_73_1_R0_clk = R0_clk;
  assign mem_73_1_R0_en = R0_en & R0_addr_sel == 8'h49;
  assign mem_73_1_W0_addr = W0_addr[25:0];
  assign mem_73_1_W0_clk = W0_clk;
  assign mem_73_1_W0_data = W0_data[15:8];
  assign mem_73_1_W0_en = W0_en & W0_addr_sel == 8'h49;
  assign mem_73_1_W0_mask = W0_mask[1];
  assign mem_73_2_R0_addr = R0_addr[25:0];
  assign mem_73_2_R0_clk = R0_clk;
  assign mem_73_2_R0_en = R0_en & R0_addr_sel == 8'h49;
  assign mem_73_2_W0_addr = W0_addr[25:0];
  assign mem_73_2_W0_clk = W0_clk;
  assign mem_73_2_W0_data = W0_data[23:16];
  assign mem_73_2_W0_en = W0_en & W0_addr_sel == 8'h49;
  assign mem_73_2_W0_mask = W0_mask[2];
  assign mem_73_3_R0_addr = R0_addr[25:0];
  assign mem_73_3_R0_clk = R0_clk;
  assign mem_73_3_R0_en = R0_en & R0_addr_sel == 8'h49;
  assign mem_73_3_W0_addr = W0_addr[25:0];
  assign mem_73_3_W0_clk = W0_clk;
  assign mem_73_3_W0_data = W0_data[31:24];
  assign mem_73_3_W0_en = W0_en & W0_addr_sel == 8'h49;
  assign mem_73_3_W0_mask = W0_mask[3];
  assign mem_73_4_R0_addr = R0_addr[25:0];
  assign mem_73_4_R0_clk = R0_clk;
  assign mem_73_4_R0_en = R0_en & R0_addr_sel == 8'h49;
  assign mem_73_4_W0_addr = W0_addr[25:0];
  assign mem_73_4_W0_clk = W0_clk;
  assign mem_73_4_W0_data = W0_data[39:32];
  assign mem_73_4_W0_en = W0_en & W0_addr_sel == 8'h49;
  assign mem_73_4_W0_mask = W0_mask[4];
  assign mem_73_5_R0_addr = R0_addr[25:0];
  assign mem_73_5_R0_clk = R0_clk;
  assign mem_73_5_R0_en = R0_en & R0_addr_sel == 8'h49;
  assign mem_73_5_W0_addr = W0_addr[25:0];
  assign mem_73_5_W0_clk = W0_clk;
  assign mem_73_5_W0_data = W0_data[47:40];
  assign mem_73_5_W0_en = W0_en & W0_addr_sel == 8'h49;
  assign mem_73_5_W0_mask = W0_mask[5];
  assign mem_73_6_R0_addr = R0_addr[25:0];
  assign mem_73_6_R0_clk = R0_clk;
  assign mem_73_6_R0_en = R0_en & R0_addr_sel == 8'h49;
  assign mem_73_6_W0_addr = W0_addr[25:0];
  assign mem_73_6_W0_clk = W0_clk;
  assign mem_73_6_W0_data = W0_data[55:48];
  assign mem_73_6_W0_en = W0_en & W0_addr_sel == 8'h49;
  assign mem_73_6_W0_mask = W0_mask[6];
  assign mem_73_7_R0_addr = R0_addr[25:0];
  assign mem_73_7_R0_clk = R0_clk;
  assign mem_73_7_R0_en = R0_en & R0_addr_sel == 8'h49;
  assign mem_73_7_W0_addr = W0_addr[25:0];
  assign mem_73_7_W0_clk = W0_clk;
  assign mem_73_7_W0_data = W0_data[63:56];
  assign mem_73_7_W0_en = W0_en & W0_addr_sel == 8'h49;
  assign mem_73_7_W0_mask = W0_mask[7];
  assign mem_74_0_R0_addr = R0_addr[25:0];
  assign mem_74_0_R0_clk = R0_clk;
  assign mem_74_0_R0_en = R0_en & R0_addr_sel == 8'h4a;
  assign mem_74_0_W0_addr = W0_addr[25:0];
  assign mem_74_0_W0_clk = W0_clk;
  assign mem_74_0_W0_data = W0_data[7:0];
  assign mem_74_0_W0_en = W0_en & W0_addr_sel == 8'h4a;
  assign mem_74_0_W0_mask = W0_mask[0];
  assign mem_74_1_R0_addr = R0_addr[25:0];
  assign mem_74_1_R0_clk = R0_clk;
  assign mem_74_1_R0_en = R0_en & R0_addr_sel == 8'h4a;
  assign mem_74_1_W0_addr = W0_addr[25:0];
  assign mem_74_1_W0_clk = W0_clk;
  assign mem_74_1_W0_data = W0_data[15:8];
  assign mem_74_1_W0_en = W0_en & W0_addr_sel == 8'h4a;
  assign mem_74_1_W0_mask = W0_mask[1];
  assign mem_74_2_R0_addr = R0_addr[25:0];
  assign mem_74_2_R0_clk = R0_clk;
  assign mem_74_2_R0_en = R0_en & R0_addr_sel == 8'h4a;
  assign mem_74_2_W0_addr = W0_addr[25:0];
  assign mem_74_2_W0_clk = W0_clk;
  assign mem_74_2_W0_data = W0_data[23:16];
  assign mem_74_2_W0_en = W0_en & W0_addr_sel == 8'h4a;
  assign mem_74_2_W0_mask = W0_mask[2];
  assign mem_74_3_R0_addr = R0_addr[25:0];
  assign mem_74_3_R0_clk = R0_clk;
  assign mem_74_3_R0_en = R0_en & R0_addr_sel == 8'h4a;
  assign mem_74_3_W0_addr = W0_addr[25:0];
  assign mem_74_3_W0_clk = W0_clk;
  assign mem_74_3_W0_data = W0_data[31:24];
  assign mem_74_3_W0_en = W0_en & W0_addr_sel == 8'h4a;
  assign mem_74_3_W0_mask = W0_mask[3];
  assign mem_74_4_R0_addr = R0_addr[25:0];
  assign mem_74_4_R0_clk = R0_clk;
  assign mem_74_4_R0_en = R0_en & R0_addr_sel == 8'h4a;
  assign mem_74_4_W0_addr = W0_addr[25:0];
  assign mem_74_4_W0_clk = W0_clk;
  assign mem_74_4_W0_data = W0_data[39:32];
  assign mem_74_4_W0_en = W0_en & W0_addr_sel == 8'h4a;
  assign mem_74_4_W0_mask = W0_mask[4];
  assign mem_74_5_R0_addr = R0_addr[25:0];
  assign mem_74_5_R0_clk = R0_clk;
  assign mem_74_5_R0_en = R0_en & R0_addr_sel == 8'h4a;
  assign mem_74_5_W0_addr = W0_addr[25:0];
  assign mem_74_5_W0_clk = W0_clk;
  assign mem_74_5_W0_data = W0_data[47:40];
  assign mem_74_5_W0_en = W0_en & W0_addr_sel == 8'h4a;
  assign mem_74_5_W0_mask = W0_mask[5];
  assign mem_74_6_R0_addr = R0_addr[25:0];
  assign mem_74_6_R0_clk = R0_clk;
  assign mem_74_6_R0_en = R0_en & R0_addr_sel == 8'h4a;
  assign mem_74_6_W0_addr = W0_addr[25:0];
  assign mem_74_6_W0_clk = W0_clk;
  assign mem_74_6_W0_data = W0_data[55:48];
  assign mem_74_6_W0_en = W0_en & W0_addr_sel == 8'h4a;
  assign mem_74_6_W0_mask = W0_mask[6];
  assign mem_74_7_R0_addr = R0_addr[25:0];
  assign mem_74_7_R0_clk = R0_clk;
  assign mem_74_7_R0_en = R0_en & R0_addr_sel == 8'h4a;
  assign mem_74_7_W0_addr = W0_addr[25:0];
  assign mem_74_7_W0_clk = W0_clk;
  assign mem_74_7_W0_data = W0_data[63:56];
  assign mem_74_7_W0_en = W0_en & W0_addr_sel == 8'h4a;
  assign mem_74_7_W0_mask = W0_mask[7];
  assign mem_75_0_R0_addr = R0_addr[25:0];
  assign mem_75_0_R0_clk = R0_clk;
  assign mem_75_0_R0_en = R0_en & R0_addr_sel == 8'h4b;
  assign mem_75_0_W0_addr = W0_addr[25:0];
  assign mem_75_0_W0_clk = W0_clk;
  assign mem_75_0_W0_data = W0_data[7:0];
  assign mem_75_0_W0_en = W0_en & W0_addr_sel == 8'h4b;
  assign mem_75_0_W0_mask = W0_mask[0];
  assign mem_75_1_R0_addr = R0_addr[25:0];
  assign mem_75_1_R0_clk = R0_clk;
  assign mem_75_1_R0_en = R0_en & R0_addr_sel == 8'h4b;
  assign mem_75_1_W0_addr = W0_addr[25:0];
  assign mem_75_1_W0_clk = W0_clk;
  assign mem_75_1_W0_data = W0_data[15:8];
  assign mem_75_1_W0_en = W0_en & W0_addr_sel == 8'h4b;
  assign mem_75_1_W0_mask = W0_mask[1];
  assign mem_75_2_R0_addr = R0_addr[25:0];
  assign mem_75_2_R0_clk = R0_clk;
  assign mem_75_2_R0_en = R0_en & R0_addr_sel == 8'h4b;
  assign mem_75_2_W0_addr = W0_addr[25:0];
  assign mem_75_2_W0_clk = W0_clk;
  assign mem_75_2_W0_data = W0_data[23:16];
  assign mem_75_2_W0_en = W0_en & W0_addr_sel == 8'h4b;
  assign mem_75_2_W0_mask = W0_mask[2];
  assign mem_75_3_R0_addr = R0_addr[25:0];
  assign mem_75_3_R0_clk = R0_clk;
  assign mem_75_3_R0_en = R0_en & R0_addr_sel == 8'h4b;
  assign mem_75_3_W0_addr = W0_addr[25:0];
  assign mem_75_3_W0_clk = W0_clk;
  assign mem_75_3_W0_data = W0_data[31:24];
  assign mem_75_3_W0_en = W0_en & W0_addr_sel == 8'h4b;
  assign mem_75_3_W0_mask = W0_mask[3];
  assign mem_75_4_R0_addr = R0_addr[25:0];
  assign mem_75_4_R0_clk = R0_clk;
  assign mem_75_4_R0_en = R0_en & R0_addr_sel == 8'h4b;
  assign mem_75_4_W0_addr = W0_addr[25:0];
  assign mem_75_4_W0_clk = W0_clk;
  assign mem_75_4_W0_data = W0_data[39:32];
  assign mem_75_4_W0_en = W0_en & W0_addr_sel == 8'h4b;
  assign mem_75_4_W0_mask = W0_mask[4];
  assign mem_75_5_R0_addr = R0_addr[25:0];
  assign mem_75_5_R0_clk = R0_clk;
  assign mem_75_5_R0_en = R0_en & R0_addr_sel == 8'h4b;
  assign mem_75_5_W0_addr = W0_addr[25:0];
  assign mem_75_5_W0_clk = W0_clk;
  assign mem_75_5_W0_data = W0_data[47:40];
  assign mem_75_5_W0_en = W0_en & W0_addr_sel == 8'h4b;
  assign mem_75_5_W0_mask = W0_mask[5];
  assign mem_75_6_R0_addr = R0_addr[25:0];
  assign mem_75_6_R0_clk = R0_clk;
  assign mem_75_6_R0_en = R0_en & R0_addr_sel == 8'h4b;
  assign mem_75_6_W0_addr = W0_addr[25:0];
  assign mem_75_6_W0_clk = W0_clk;
  assign mem_75_6_W0_data = W0_data[55:48];
  assign mem_75_6_W0_en = W0_en & W0_addr_sel == 8'h4b;
  assign mem_75_6_W0_mask = W0_mask[6];
  assign mem_75_7_R0_addr = R0_addr[25:0];
  assign mem_75_7_R0_clk = R0_clk;
  assign mem_75_7_R0_en = R0_en & R0_addr_sel == 8'h4b;
  assign mem_75_7_W0_addr = W0_addr[25:0];
  assign mem_75_7_W0_clk = W0_clk;
  assign mem_75_7_W0_data = W0_data[63:56];
  assign mem_75_7_W0_en = W0_en & W0_addr_sel == 8'h4b;
  assign mem_75_7_W0_mask = W0_mask[7];
  assign mem_76_0_R0_addr = R0_addr[25:0];
  assign mem_76_0_R0_clk = R0_clk;
  assign mem_76_0_R0_en = R0_en & R0_addr_sel == 8'h4c;
  assign mem_76_0_W0_addr = W0_addr[25:0];
  assign mem_76_0_W0_clk = W0_clk;
  assign mem_76_0_W0_data = W0_data[7:0];
  assign mem_76_0_W0_en = W0_en & W0_addr_sel == 8'h4c;
  assign mem_76_0_W0_mask = W0_mask[0];
  assign mem_76_1_R0_addr = R0_addr[25:0];
  assign mem_76_1_R0_clk = R0_clk;
  assign mem_76_1_R0_en = R0_en & R0_addr_sel == 8'h4c;
  assign mem_76_1_W0_addr = W0_addr[25:0];
  assign mem_76_1_W0_clk = W0_clk;
  assign mem_76_1_W0_data = W0_data[15:8];
  assign mem_76_1_W0_en = W0_en & W0_addr_sel == 8'h4c;
  assign mem_76_1_W0_mask = W0_mask[1];
  assign mem_76_2_R0_addr = R0_addr[25:0];
  assign mem_76_2_R0_clk = R0_clk;
  assign mem_76_2_R0_en = R0_en & R0_addr_sel == 8'h4c;
  assign mem_76_2_W0_addr = W0_addr[25:0];
  assign mem_76_2_W0_clk = W0_clk;
  assign mem_76_2_W0_data = W0_data[23:16];
  assign mem_76_2_W0_en = W0_en & W0_addr_sel == 8'h4c;
  assign mem_76_2_W0_mask = W0_mask[2];
  assign mem_76_3_R0_addr = R0_addr[25:0];
  assign mem_76_3_R0_clk = R0_clk;
  assign mem_76_3_R0_en = R0_en & R0_addr_sel == 8'h4c;
  assign mem_76_3_W0_addr = W0_addr[25:0];
  assign mem_76_3_W0_clk = W0_clk;
  assign mem_76_3_W0_data = W0_data[31:24];
  assign mem_76_3_W0_en = W0_en & W0_addr_sel == 8'h4c;
  assign mem_76_3_W0_mask = W0_mask[3];
  assign mem_76_4_R0_addr = R0_addr[25:0];
  assign mem_76_4_R0_clk = R0_clk;
  assign mem_76_4_R0_en = R0_en & R0_addr_sel == 8'h4c;
  assign mem_76_4_W0_addr = W0_addr[25:0];
  assign mem_76_4_W0_clk = W0_clk;
  assign mem_76_4_W0_data = W0_data[39:32];
  assign mem_76_4_W0_en = W0_en & W0_addr_sel == 8'h4c;
  assign mem_76_4_W0_mask = W0_mask[4];
  assign mem_76_5_R0_addr = R0_addr[25:0];
  assign mem_76_5_R0_clk = R0_clk;
  assign mem_76_5_R0_en = R0_en & R0_addr_sel == 8'h4c;
  assign mem_76_5_W0_addr = W0_addr[25:0];
  assign mem_76_5_W0_clk = W0_clk;
  assign mem_76_5_W0_data = W0_data[47:40];
  assign mem_76_5_W0_en = W0_en & W0_addr_sel == 8'h4c;
  assign mem_76_5_W0_mask = W0_mask[5];
  assign mem_76_6_R0_addr = R0_addr[25:0];
  assign mem_76_6_R0_clk = R0_clk;
  assign mem_76_6_R0_en = R0_en & R0_addr_sel == 8'h4c;
  assign mem_76_6_W0_addr = W0_addr[25:0];
  assign mem_76_6_W0_clk = W0_clk;
  assign mem_76_6_W0_data = W0_data[55:48];
  assign mem_76_6_W0_en = W0_en & W0_addr_sel == 8'h4c;
  assign mem_76_6_W0_mask = W0_mask[6];
  assign mem_76_7_R0_addr = R0_addr[25:0];
  assign mem_76_7_R0_clk = R0_clk;
  assign mem_76_7_R0_en = R0_en & R0_addr_sel == 8'h4c;
  assign mem_76_7_W0_addr = W0_addr[25:0];
  assign mem_76_7_W0_clk = W0_clk;
  assign mem_76_7_W0_data = W0_data[63:56];
  assign mem_76_7_W0_en = W0_en & W0_addr_sel == 8'h4c;
  assign mem_76_7_W0_mask = W0_mask[7];
  assign mem_77_0_R0_addr = R0_addr[25:0];
  assign mem_77_0_R0_clk = R0_clk;
  assign mem_77_0_R0_en = R0_en & R0_addr_sel == 8'h4d;
  assign mem_77_0_W0_addr = W0_addr[25:0];
  assign mem_77_0_W0_clk = W0_clk;
  assign mem_77_0_W0_data = W0_data[7:0];
  assign mem_77_0_W0_en = W0_en & W0_addr_sel == 8'h4d;
  assign mem_77_0_W0_mask = W0_mask[0];
  assign mem_77_1_R0_addr = R0_addr[25:0];
  assign mem_77_1_R0_clk = R0_clk;
  assign mem_77_1_R0_en = R0_en & R0_addr_sel == 8'h4d;
  assign mem_77_1_W0_addr = W0_addr[25:0];
  assign mem_77_1_W0_clk = W0_clk;
  assign mem_77_1_W0_data = W0_data[15:8];
  assign mem_77_1_W0_en = W0_en & W0_addr_sel == 8'h4d;
  assign mem_77_1_W0_mask = W0_mask[1];
  assign mem_77_2_R0_addr = R0_addr[25:0];
  assign mem_77_2_R0_clk = R0_clk;
  assign mem_77_2_R0_en = R0_en & R0_addr_sel == 8'h4d;
  assign mem_77_2_W0_addr = W0_addr[25:0];
  assign mem_77_2_W0_clk = W0_clk;
  assign mem_77_2_W0_data = W0_data[23:16];
  assign mem_77_2_W0_en = W0_en & W0_addr_sel == 8'h4d;
  assign mem_77_2_W0_mask = W0_mask[2];
  assign mem_77_3_R0_addr = R0_addr[25:0];
  assign mem_77_3_R0_clk = R0_clk;
  assign mem_77_3_R0_en = R0_en & R0_addr_sel == 8'h4d;
  assign mem_77_3_W0_addr = W0_addr[25:0];
  assign mem_77_3_W0_clk = W0_clk;
  assign mem_77_3_W0_data = W0_data[31:24];
  assign mem_77_3_W0_en = W0_en & W0_addr_sel == 8'h4d;
  assign mem_77_3_W0_mask = W0_mask[3];
  assign mem_77_4_R0_addr = R0_addr[25:0];
  assign mem_77_4_R0_clk = R0_clk;
  assign mem_77_4_R0_en = R0_en & R0_addr_sel == 8'h4d;
  assign mem_77_4_W0_addr = W0_addr[25:0];
  assign mem_77_4_W0_clk = W0_clk;
  assign mem_77_4_W0_data = W0_data[39:32];
  assign mem_77_4_W0_en = W0_en & W0_addr_sel == 8'h4d;
  assign mem_77_4_W0_mask = W0_mask[4];
  assign mem_77_5_R0_addr = R0_addr[25:0];
  assign mem_77_5_R0_clk = R0_clk;
  assign mem_77_5_R0_en = R0_en & R0_addr_sel == 8'h4d;
  assign mem_77_5_W0_addr = W0_addr[25:0];
  assign mem_77_5_W0_clk = W0_clk;
  assign mem_77_5_W0_data = W0_data[47:40];
  assign mem_77_5_W0_en = W0_en & W0_addr_sel == 8'h4d;
  assign mem_77_5_W0_mask = W0_mask[5];
  assign mem_77_6_R0_addr = R0_addr[25:0];
  assign mem_77_6_R0_clk = R0_clk;
  assign mem_77_6_R0_en = R0_en & R0_addr_sel == 8'h4d;
  assign mem_77_6_W0_addr = W0_addr[25:0];
  assign mem_77_6_W0_clk = W0_clk;
  assign mem_77_6_W0_data = W0_data[55:48];
  assign mem_77_6_W0_en = W0_en & W0_addr_sel == 8'h4d;
  assign mem_77_6_W0_mask = W0_mask[6];
  assign mem_77_7_R0_addr = R0_addr[25:0];
  assign mem_77_7_R0_clk = R0_clk;
  assign mem_77_7_R0_en = R0_en & R0_addr_sel == 8'h4d;
  assign mem_77_7_W0_addr = W0_addr[25:0];
  assign mem_77_7_W0_clk = W0_clk;
  assign mem_77_7_W0_data = W0_data[63:56];
  assign mem_77_7_W0_en = W0_en & W0_addr_sel == 8'h4d;
  assign mem_77_7_W0_mask = W0_mask[7];
  assign mem_78_0_R0_addr = R0_addr[25:0];
  assign mem_78_0_R0_clk = R0_clk;
  assign mem_78_0_R0_en = R0_en & R0_addr_sel == 8'h4e;
  assign mem_78_0_W0_addr = W0_addr[25:0];
  assign mem_78_0_W0_clk = W0_clk;
  assign mem_78_0_W0_data = W0_data[7:0];
  assign mem_78_0_W0_en = W0_en & W0_addr_sel == 8'h4e;
  assign mem_78_0_W0_mask = W0_mask[0];
  assign mem_78_1_R0_addr = R0_addr[25:0];
  assign mem_78_1_R0_clk = R0_clk;
  assign mem_78_1_R0_en = R0_en & R0_addr_sel == 8'h4e;
  assign mem_78_1_W0_addr = W0_addr[25:0];
  assign mem_78_1_W0_clk = W0_clk;
  assign mem_78_1_W0_data = W0_data[15:8];
  assign mem_78_1_W0_en = W0_en & W0_addr_sel == 8'h4e;
  assign mem_78_1_W0_mask = W0_mask[1];
  assign mem_78_2_R0_addr = R0_addr[25:0];
  assign mem_78_2_R0_clk = R0_clk;
  assign mem_78_2_R0_en = R0_en & R0_addr_sel == 8'h4e;
  assign mem_78_2_W0_addr = W0_addr[25:0];
  assign mem_78_2_W0_clk = W0_clk;
  assign mem_78_2_W0_data = W0_data[23:16];
  assign mem_78_2_W0_en = W0_en & W0_addr_sel == 8'h4e;
  assign mem_78_2_W0_mask = W0_mask[2];
  assign mem_78_3_R0_addr = R0_addr[25:0];
  assign mem_78_3_R0_clk = R0_clk;
  assign mem_78_3_R0_en = R0_en & R0_addr_sel == 8'h4e;
  assign mem_78_3_W0_addr = W0_addr[25:0];
  assign mem_78_3_W0_clk = W0_clk;
  assign mem_78_3_W0_data = W0_data[31:24];
  assign mem_78_3_W0_en = W0_en & W0_addr_sel == 8'h4e;
  assign mem_78_3_W0_mask = W0_mask[3];
  assign mem_78_4_R0_addr = R0_addr[25:0];
  assign mem_78_4_R0_clk = R0_clk;
  assign mem_78_4_R0_en = R0_en & R0_addr_sel == 8'h4e;
  assign mem_78_4_W0_addr = W0_addr[25:0];
  assign mem_78_4_W0_clk = W0_clk;
  assign mem_78_4_W0_data = W0_data[39:32];
  assign mem_78_4_W0_en = W0_en & W0_addr_sel == 8'h4e;
  assign mem_78_4_W0_mask = W0_mask[4];
  assign mem_78_5_R0_addr = R0_addr[25:0];
  assign mem_78_5_R0_clk = R0_clk;
  assign mem_78_5_R0_en = R0_en & R0_addr_sel == 8'h4e;
  assign mem_78_5_W0_addr = W0_addr[25:0];
  assign mem_78_5_W0_clk = W0_clk;
  assign mem_78_5_W0_data = W0_data[47:40];
  assign mem_78_5_W0_en = W0_en & W0_addr_sel == 8'h4e;
  assign mem_78_5_W0_mask = W0_mask[5];
  assign mem_78_6_R0_addr = R0_addr[25:0];
  assign mem_78_6_R0_clk = R0_clk;
  assign mem_78_6_R0_en = R0_en & R0_addr_sel == 8'h4e;
  assign mem_78_6_W0_addr = W0_addr[25:0];
  assign mem_78_6_W0_clk = W0_clk;
  assign mem_78_6_W0_data = W0_data[55:48];
  assign mem_78_6_W0_en = W0_en & W0_addr_sel == 8'h4e;
  assign mem_78_6_W0_mask = W0_mask[6];
  assign mem_78_7_R0_addr = R0_addr[25:0];
  assign mem_78_7_R0_clk = R0_clk;
  assign mem_78_7_R0_en = R0_en & R0_addr_sel == 8'h4e;
  assign mem_78_7_W0_addr = W0_addr[25:0];
  assign mem_78_7_W0_clk = W0_clk;
  assign mem_78_7_W0_data = W0_data[63:56];
  assign mem_78_7_W0_en = W0_en & W0_addr_sel == 8'h4e;
  assign mem_78_7_W0_mask = W0_mask[7];
  assign mem_79_0_R0_addr = R0_addr[25:0];
  assign mem_79_0_R0_clk = R0_clk;
  assign mem_79_0_R0_en = R0_en & R0_addr_sel == 8'h4f;
  assign mem_79_0_W0_addr = W0_addr[25:0];
  assign mem_79_0_W0_clk = W0_clk;
  assign mem_79_0_W0_data = W0_data[7:0];
  assign mem_79_0_W0_en = W0_en & W0_addr_sel == 8'h4f;
  assign mem_79_0_W0_mask = W0_mask[0];
  assign mem_79_1_R0_addr = R0_addr[25:0];
  assign mem_79_1_R0_clk = R0_clk;
  assign mem_79_1_R0_en = R0_en & R0_addr_sel == 8'h4f;
  assign mem_79_1_W0_addr = W0_addr[25:0];
  assign mem_79_1_W0_clk = W0_clk;
  assign mem_79_1_W0_data = W0_data[15:8];
  assign mem_79_1_W0_en = W0_en & W0_addr_sel == 8'h4f;
  assign mem_79_1_W0_mask = W0_mask[1];
  assign mem_79_2_R0_addr = R0_addr[25:0];
  assign mem_79_2_R0_clk = R0_clk;
  assign mem_79_2_R0_en = R0_en & R0_addr_sel == 8'h4f;
  assign mem_79_2_W0_addr = W0_addr[25:0];
  assign mem_79_2_W0_clk = W0_clk;
  assign mem_79_2_W0_data = W0_data[23:16];
  assign mem_79_2_W0_en = W0_en & W0_addr_sel == 8'h4f;
  assign mem_79_2_W0_mask = W0_mask[2];
  assign mem_79_3_R0_addr = R0_addr[25:0];
  assign mem_79_3_R0_clk = R0_clk;
  assign mem_79_3_R0_en = R0_en & R0_addr_sel == 8'h4f;
  assign mem_79_3_W0_addr = W0_addr[25:0];
  assign mem_79_3_W0_clk = W0_clk;
  assign mem_79_3_W0_data = W0_data[31:24];
  assign mem_79_3_W0_en = W0_en & W0_addr_sel == 8'h4f;
  assign mem_79_3_W0_mask = W0_mask[3];
  assign mem_79_4_R0_addr = R0_addr[25:0];
  assign mem_79_4_R0_clk = R0_clk;
  assign mem_79_4_R0_en = R0_en & R0_addr_sel == 8'h4f;
  assign mem_79_4_W0_addr = W0_addr[25:0];
  assign mem_79_4_W0_clk = W0_clk;
  assign mem_79_4_W0_data = W0_data[39:32];
  assign mem_79_4_W0_en = W0_en & W0_addr_sel == 8'h4f;
  assign mem_79_4_W0_mask = W0_mask[4];
  assign mem_79_5_R0_addr = R0_addr[25:0];
  assign mem_79_5_R0_clk = R0_clk;
  assign mem_79_5_R0_en = R0_en & R0_addr_sel == 8'h4f;
  assign mem_79_5_W0_addr = W0_addr[25:0];
  assign mem_79_5_W0_clk = W0_clk;
  assign mem_79_5_W0_data = W0_data[47:40];
  assign mem_79_5_W0_en = W0_en & W0_addr_sel == 8'h4f;
  assign mem_79_5_W0_mask = W0_mask[5];
  assign mem_79_6_R0_addr = R0_addr[25:0];
  assign mem_79_6_R0_clk = R0_clk;
  assign mem_79_6_R0_en = R0_en & R0_addr_sel == 8'h4f;
  assign mem_79_6_W0_addr = W0_addr[25:0];
  assign mem_79_6_W0_clk = W0_clk;
  assign mem_79_6_W0_data = W0_data[55:48];
  assign mem_79_6_W0_en = W0_en & W0_addr_sel == 8'h4f;
  assign mem_79_6_W0_mask = W0_mask[6];
  assign mem_79_7_R0_addr = R0_addr[25:0];
  assign mem_79_7_R0_clk = R0_clk;
  assign mem_79_7_R0_en = R0_en & R0_addr_sel == 8'h4f;
  assign mem_79_7_W0_addr = W0_addr[25:0];
  assign mem_79_7_W0_clk = W0_clk;
  assign mem_79_7_W0_data = W0_data[63:56];
  assign mem_79_7_W0_en = W0_en & W0_addr_sel == 8'h4f;
  assign mem_79_7_W0_mask = W0_mask[7];
  assign mem_80_0_R0_addr = R0_addr[25:0];
  assign mem_80_0_R0_clk = R0_clk;
  assign mem_80_0_R0_en = R0_en & R0_addr_sel == 8'h50;
  assign mem_80_0_W0_addr = W0_addr[25:0];
  assign mem_80_0_W0_clk = W0_clk;
  assign mem_80_0_W0_data = W0_data[7:0];
  assign mem_80_0_W0_en = W0_en & W0_addr_sel == 8'h50;
  assign mem_80_0_W0_mask = W0_mask[0];
  assign mem_80_1_R0_addr = R0_addr[25:0];
  assign mem_80_1_R0_clk = R0_clk;
  assign mem_80_1_R0_en = R0_en & R0_addr_sel == 8'h50;
  assign mem_80_1_W0_addr = W0_addr[25:0];
  assign mem_80_1_W0_clk = W0_clk;
  assign mem_80_1_W0_data = W0_data[15:8];
  assign mem_80_1_W0_en = W0_en & W0_addr_sel == 8'h50;
  assign mem_80_1_W0_mask = W0_mask[1];
  assign mem_80_2_R0_addr = R0_addr[25:0];
  assign mem_80_2_R0_clk = R0_clk;
  assign mem_80_2_R0_en = R0_en & R0_addr_sel == 8'h50;
  assign mem_80_2_W0_addr = W0_addr[25:0];
  assign mem_80_2_W0_clk = W0_clk;
  assign mem_80_2_W0_data = W0_data[23:16];
  assign mem_80_2_W0_en = W0_en & W0_addr_sel == 8'h50;
  assign mem_80_2_W0_mask = W0_mask[2];
  assign mem_80_3_R0_addr = R0_addr[25:0];
  assign mem_80_3_R0_clk = R0_clk;
  assign mem_80_3_R0_en = R0_en & R0_addr_sel == 8'h50;
  assign mem_80_3_W0_addr = W0_addr[25:0];
  assign mem_80_3_W0_clk = W0_clk;
  assign mem_80_3_W0_data = W0_data[31:24];
  assign mem_80_3_W0_en = W0_en & W0_addr_sel == 8'h50;
  assign mem_80_3_W0_mask = W0_mask[3];
  assign mem_80_4_R0_addr = R0_addr[25:0];
  assign mem_80_4_R0_clk = R0_clk;
  assign mem_80_4_R0_en = R0_en & R0_addr_sel == 8'h50;
  assign mem_80_4_W0_addr = W0_addr[25:0];
  assign mem_80_4_W0_clk = W0_clk;
  assign mem_80_4_W0_data = W0_data[39:32];
  assign mem_80_4_W0_en = W0_en & W0_addr_sel == 8'h50;
  assign mem_80_4_W0_mask = W0_mask[4];
  assign mem_80_5_R0_addr = R0_addr[25:0];
  assign mem_80_5_R0_clk = R0_clk;
  assign mem_80_5_R0_en = R0_en & R0_addr_sel == 8'h50;
  assign mem_80_5_W0_addr = W0_addr[25:0];
  assign mem_80_5_W0_clk = W0_clk;
  assign mem_80_5_W0_data = W0_data[47:40];
  assign mem_80_5_W0_en = W0_en & W0_addr_sel == 8'h50;
  assign mem_80_5_W0_mask = W0_mask[5];
  assign mem_80_6_R0_addr = R0_addr[25:0];
  assign mem_80_6_R0_clk = R0_clk;
  assign mem_80_6_R0_en = R0_en & R0_addr_sel == 8'h50;
  assign mem_80_6_W0_addr = W0_addr[25:0];
  assign mem_80_6_W0_clk = W0_clk;
  assign mem_80_6_W0_data = W0_data[55:48];
  assign mem_80_6_W0_en = W0_en & W0_addr_sel == 8'h50;
  assign mem_80_6_W0_mask = W0_mask[6];
  assign mem_80_7_R0_addr = R0_addr[25:0];
  assign mem_80_7_R0_clk = R0_clk;
  assign mem_80_7_R0_en = R0_en & R0_addr_sel == 8'h50;
  assign mem_80_7_W0_addr = W0_addr[25:0];
  assign mem_80_7_W0_clk = W0_clk;
  assign mem_80_7_W0_data = W0_data[63:56];
  assign mem_80_7_W0_en = W0_en & W0_addr_sel == 8'h50;
  assign mem_80_7_W0_mask = W0_mask[7];
  assign mem_81_0_R0_addr = R0_addr[25:0];
  assign mem_81_0_R0_clk = R0_clk;
  assign mem_81_0_R0_en = R0_en & R0_addr_sel == 8'h51;
  assign mem_81_0_W0_addr = W0_addr[25:0];
  assign mem_81_0_W0_clk = W0_clk;
  assign mem_81_0_W0_data = W0_data[7:0];
  assign mem_81_0_W0_en = W0_en & W0_addr_sel == 8'h51;
  assign mem_81_0_W0_mask = W0_mask[0];
  assign mem_81_1_R0_addr = R0_addr[25:0];
  assign mem_81_1_R0_clk = R0_clk;
  assign mem_81_1_R0_en = R0_en & R0_addr_sel == 8'h51;
  assign mem_81_1_W0_addr = W0_addr[25:0];
  assign mem_81_1_W0_clk = W0_clk;
  assign mem_81_1_W0_data = W0_data[15:8];
  assign mem_81_1_W0_en = W0_en & W0_addr_sel == 8'h51;
  assign mem_81_1_W0_mask = W0_mask[1];
  assign mem_81_2_R0_addr = R0_addr[25:0];
  assign mem_81_2_R0_clk = R0_clk;
  assign mem_81_2_R0_en = R0_en & R0_addr_sel == 8'h51;
  assign mem_81_2_W0_addr = W0_addr[25:0];
  assign mem_81_2_W0_clk = W0_clk;
  assign mem_81_2_W0_data = W0_data[23:16];
  assign mem_81_2_W0_en = W0_en & W0_addr_sel == 8'h51;
  assign mem_81_2_W0_mask = W0_mask[2];
  assign mem_81_3_R0_addr = R0_addr[25:0];
  assign mem_81_3_R0_clk = R0_clk;
  assign mem_81_3_R0_en = R0_en & R0_addr_sel == 8'h51;
  assign mem_81_3_W0_addr = W0_addr[25:0];
  assign mem_81_3_W0_clk = W0_clk;
  assign mem_81_3_W0_data = W0_data[31:24];
  assign mem_81_3_W0_en = W0_en & W0_addr_sel == 8'h51;
  assign mem_81_3_W0_mask = W0_mask[3];
  assign mem_81_4_R0_addr = R0_addr[25:0];
  assign mem_81_4_R0_clk = R0_clk;
  assign mem_81_4_R0_en = R0_en & R0_addr_sel == 8'h51;
  assign mem_81_4_W0_addr = W0_addr[25:0];
  assign mem_81_4_W0_clk = W0_clk;
  assign mem_81_4_W0_data = W0_data[39:32];
  assign mem_81_4_W0_en = W0_en & W0_addr_sel == 8'h51;
  assign mem_81_4_W0_mask = W0_mask[4];
  assign mem_81_5_R0_addr = R0_addr[25:0];
  assign mem_81_5_R0_clk = R0_clk;
  assign mem_81_5_R0_en = R0_en & R0_addr_sel == 8'h51;
  assign mem_81_5_W0_addr = W0_addr[25:0];
  assign mem_81_5_W0_clk = W0_clk;
  assign mem_81_5_W0_data = W0_data[47:40];
  assign mem_81_5_W0_en = W0_en & W0_addr_sel == 8'h51;
  assign mem_81_5_W0_mask = W0_mask[5];
  assign mem_81_6_R0_addr = R0_addr[25:0];
  assign mem_81_6_R0_clk = R0_clk;
  assign mem_81_6_R0_en = R0_en & R0_addr_sel == 8'h51;
  assign mem_81_6_W0_addr = W0_addr[25:0];
  assign mem_81_6_W0_clk = W0_clk;
  assign mem_81_6_W0_data = W0_data[55:48];
  assign mem_81_6_W0_en = W0_en & W0_addr_sel == 8'h51;
  assign mem_81_6_W0_mask = W0_mask[6];
  assign mem_81_7_R0_addr = R0_addr[25:0];
  assign mem_81_7_R0_clk = R0_clk;
  assign mem_81_7_R0_en = R0_en & R0_addr_sel == 8'h51;
  assign mem_81_7_W0_addr = W0_addr[25:0];
  assign mem_81_7_W0_clk = W0_clk;
  assign mem_81_7_W0_data = W0_data[63:56];
  assign mem_81_7_W0_en = W0_en & W0_addr_sel == 8'h51;
  assign mem_81_7_W0_mask = W0_mask[7];
  assign mem_82_0_R0_addr = R0_addr[25:0];
  assign mem_82_0_R0_clk = R0_clk;
  assign mem_82_0_R0_en = R0_en & R0_addr_sel == 8'h52;
  assign mem_82_0_W0_addr = W0_addr[25:0];
  assign mem_82_0_W0_clk = W0_clk;
  assign mem_82_0_W0_data = W0_data[7:0];
  assign mem_82_0_W0_en = W0_en & W0_addr_sel == 8'h52;
  assign mem_82_0_W0_mask = W0_mask[0];
  assign mem_82_1_R0_addr = R0_addr[25:0];
  assign mem_82_1_R0_clk = R0_clk;
  assign mem_82_1_R0_en = R0_en & R0_addr_sel == 8'h52;
  assign mem_82_1_W0_addr = W0_addr[25:0];
  assign mem_82_1_W0_clk = W0_clk;
  assign mem_82_1_W0_data = W0_data[15:8];
  assign mem_82_1_W0_en = W0_en & W0_addr_sel == 8'h52;
  assign mem_82_1_W0_mask = W0_mask[1];
  assign mem_82_2_R0_addr = R0_addr[25:0];
  assign mem_82_2_R0_clk = R0_clk;
  assign mem_82_2_R0_en = R0_en & R0_addr_sel == 8'h52;
  assign mem_82_2_W0_addr = W0_addr[25:0];
  assign mem_82_2_W0_clk = W0_clk;
  assign mem_82_2_W0_data = W0_data[23:16];
  assign mem_82_2_W0_en = W0_en & W0_addr_sel == 8'h52;
  assign mem_82_2_W0_mask = W0_mask[2];
  assign mem_82_3_R0_addr = R0_addr[25:0];
  assign mem_82_3_R0_clk = R0_clk;
  assign mem_82_3_R0_en = R0_en & R0_addr_sel == 8'h52;
  assign mem_82_3_W0_addr = W0_addr[25:0];
  assign mem_82_3_W0_clk = W0_clk;
  assign mem_82_3_W0_data = W0_data[31:24];
  assign mem_82_3_W0_en = W0_en & W0_addr_sel == 8'h52;
  assign mem_82_3_W0_mask = W0_mask[3];
  assign mem_82_4_R0_addr = R0_addr[25:0];
  assign mem_82_4_R0_clk = R0_clk;
  assign mem_82_4_R0_en = R0_en & R0_addr_sel == 8'h52;
  assign mem_82_4_W0_addr = W0_addr[25:0];
  assign mem_82_4_W0_clk = W0_clk;
  assign mem_82_4_W0_data = W0_data[39:32];
  assign mem_82_4_W0_en = W0_en & W0_addr_sel == 8'h52;
  assign mem_82_4_W0_mask = W0_mask[4];
  assign mem_82_5_R0_addr = R0_addr[25:0];
  assign mem_82_5_R0_clk = R0_clk;
  assign mem_82_5_R0_en = R0_en & R0_addr_sel == 8'h52;
  assign mem_82_5_W0_addr = W0_addr[25:0];
  assign mem_82_5_W0_clk = W0_clk;
  assign mem_82_5_W0_data = W0_data[47:40];
  assign mem_82_5_W0_en = W0_en & W0_addr_sel == 8'h52;
  assign mem_82_5_W0_mask = W0_mask[5];
  assign mem_82_6_R0_addr = R0_addr[25:0];
  assign mem_82_6_R0_clk = R0_clk;
  assign mem_82_6_R0_en = R0_en & R0_addr_sel == 8'h52;
  assign mem_82_6_W0_addr = W0_addr[25:0];
  assign mem_82_6_W0_clk = W0_clk;
  assign mem_82_6_W0_data = W0_data[55:48];
  assign mem_82_6_W0_en = W0_en & W0_addr_sel == 8'h52;
  assign mem_82_6_W0_mask = W0_mask[6];
  assign mem_82_7_R0_addr = R0_addr[25:0];
  assign mem_82_7_R0_clk = R0_clk;
  assign mem_82_7_R0_en = R0_en & R0_addr_sel == 8'h52;
  assign mem_82_7_W0_addr = W0_addr[25:0];
  assign mem_82_7_W0_clk = W0_clk;
  assign mem_82_7_W0_data = W0_data[63:56];
  assign mem_82_7_W0_en = W0_en & W0_addr_sel == 8'h52;
  assign mem_82_7_W0_mask = W0_mask[7];
  assign mem_83_0_R0_addr = R0_addr[25:0];
  assign mem_83_0_R0_clk = R0_clk;
  assign mem_83_0_R0_en = R0_en & R0_addr_sel == 8'h53;
  assign mem_83_0_W0_addr = W0_addr[25:0];
  assign mem_83_0_W0_clk = W0_clk;
  assign mem_83_0_W0_data = W0_data[7:0];
  assign mem_83_0_W0_en = W0_en & W0_addr_sel == 8'h53;
  assign mem_83_0_W0_mask = W0_mask[0];
  assign mem_83_1_R0_addr = R0_addr[25:0];
  assign mem_83_1_R0_clk = R0_clk;
  assign mem_83_1_R0_en = R0_en & R0_addr_sel == 8'h53;
  assign mem_83_1_W0_addr = W0_addr[25:0];
  assign mem_83_1_W0_clk = W0_clk;
  assign mem_83_1_W0_data = W0_data[15:8];
  assign mem_83_1_W0_en = W0_en & W0_addr_sel == 8'h53;
  assign mem_83_1_W0_mask = W0_mask[1];
  assign mem_83_2_R0_addr = R0_addr[25:0];
  assign mem_83_2_R0_clk = R0_clk;
  assign mem_83_2_R0_en = R0_en & R0_addr_sel == 8'h53;
  assign mem_83_2_W0_addr = W0_addr[25:0];
  assign mem_83_2_W0_clk = W0_clk;
  assign mem_83_2_W0_data = W0_data[23:16];
  assign mem_83_2_W0_en = W0_en & W0_addr_sel == 8'h53;
  assign mem_83_2_W0_mask = W0_mask[2];
  assign mem_83_3_R0_addr = R0_addr[25:0];
  assign mem_83_3_R0_clk = R0_clk;
  assign mem_83_3_R0_en = R0_en & R0_addr_sel == 8'h53;
  assign mem_83_3_W0_addr = W0_addr[25:0];
  assign mem_83_3_W0_clk = W0_clk;
  assign mem_83_3_W0_data = W0_data[31:24];
  assign mem_83_3_W0_en = W0_en & W0_addr_sel == 8'h53;
  assign mem_83_3_W0_mask = W0_mask[3];
  assign mem_83_4_R0_addr = R0_addr[25:0];
  assign mem_83_4_R0_clk = R0_clk;
  assign mem_83_4_R0_en = R0_en & R0_addr_sel == 8'h53;
  assign mem_83_4_W0_addr = W0_addr[25:0];
  assign mem_83_4_W0_clk = W0_clk;
  assign mem_83_4_W0_data = W0_data[39:32];
  assign mem_83_4_W0_en = W0_en & W0_addr_sel == 8'h53;
  assign mem_83_4_W0_mask = W0_mask[4];
  assign mem_83_5_R0_addr = R0_addr[25:0];
  assign mem_83_5_R0_clk = R0_clk;
  assign mem_83_5_R0_en = R0_en & R0_addr_sel == 8'h53;
  assign mem_83_5_W0_addr = W0_addr[25:0];
  assign mem_83_5_W0_clk = W0_clk;
  assign mem_83_5_W0_data = W0_data[47:40];
  assign mem_83_5_W0_en = W0_en & W0_addr_sel == 8'h53;
  assign mem_83_5_W0_mask = W0_mask[5];
  assign mem_83_6_R0_addr = R0_addr[25:0];
  assign mem_83_6_R0_clk = R0_clk;
  assign mem_83_6_R0_en = R0_en & R0_addr_sel == 8'h53;
  assign mem_83_6_W0_addr = W0_addr[25:0];
  assign mem_83_6_W0_clk = W0_clk;
  assign mem_83_6_W0_data = W0_data[55:48];
  assign mem_83_6_W0_en = W0_en & W0_addr_sel == 8'h53;
  assign mem_83_6_W0_mask = W0_mask[6];
  assign mem_83_7_R0_addr = R0_addr[25:0];
  assign mem_83_7_R0_clk = R0_clk;
  assign mem_83_7_R0_en = R0_en & R0_addr_sel == 8'h53;
  assign mem_83_7_W0_addr = W0_addr[25:0];
  assign mem_83_7_W0_clk = W0_clk;
  assign mem_83_7_W0_data = W0_data[63:56];
  assign mem_83_7_W0_en = W0_en & W0_addr_sel == 8'h53;
  assign mem_83_7_W0_mask = W0_mask[7];
  assign mem_84_0_R0_addr = R0_addr[25:0];
  assign mem_84_0_R0_clk = R0_clk;
  assign mem_84_0_R0_en = R0_en & R0_addr_sel == 8'h54;
  assign mem_84_0_W0_addr = W0_addr[25:0];
  assign mem_84_0_W0_clk = W0_clk;
  assign mem_84_0_W0_data = W0_data[7:0];
  assign mem_84_0_W0_en = W0_en & W0_addr_sel == 8'h54;
  assign mem_84_0_W0_mask = W0_mask[0];
  assign mem_84_1_R0_addr = R0_addr[25:0];
  assign mem_84_1_R0_clk = R0_clk;
  assign mem_84_1_R0_en = R0_en & R0_addr_sel == 8'h54;
  assign mem_84_1_W0_addr = W0_addr[25:0];
  assign mem_84_1_W0_clk = W0_clk;
  assign mem_84_1_W0_data = W0_data[15:8];
  assign mem_84_1_W0_en = W0_en & W0_addr_sel == 8'h54;
  assign mem_84_1_W0_mask = W0_mask[1];
  assign mem_84_2_R0_addr = R0_addr[25:0];
  assign mem_84_2_R0_clk = R0_clk;
  assign mem_84_2_R0_en = R0_en & R0_addr_sel == 8'h54;
  assign mem_84_2_W0_addr = W0_addr[25:0];
  assign mem_84_2_W0_clk = W0_clk;
  assign mem_84_2_W0_data = W0_data[23:16];
  assign mem_84_2_W0_en = W0_en & W0_addr_sel == 8'h54;
  assign mem_84_2_W0_mask = W0_mask[2];
  assign mem_84_3_R0_addr = R0_addr[25:0];
  assign mem_84_3_R0_clk = R0_clk;
  assign mem_84_3_R0_en = R0_en & R0_addr_sel == 8'h54;
  assign mem_84_3_W0_addr = W0_addr[25:0];
  assign mem_84_3_W0_clk = W0_clk;
  assign mem_84_3_W0_data = W0_data[31:24];
  assign mem_84_3_W0_en = W0_en & W0_addr_sel == 8'h54;
  assign mem_84_3_W0_mask = W0_mask[3];
  assign mem_84_4_R0_addr = R0_addr[25:0];
  assign mem_84_4_R0_clk = R0_clk;
  assign mem_84_4_R0_en = R0_en & R0_addr_sel == 8'h54;
  assign mem_84_4_W0_addr = W0_addr[25:0];
  assign mem_84_4_W0_clk = W0_clk;
  assign mem_84_4_W0_data = W0_data[39:32];
  assign mem_84_4_W0_en = W0_en & W0_addr_sel == 8'h54;
  assign mem_84_4_W0_mask = W0_mask[4];
  assign mem_84_5_R0_addr = R0_addr[25:0];
  assign mem_84_5_R0_clk = R0_clk;
  assign mem_84_5_R0_en = R0_en & R0_addr_sel == 8'h54;
  assign mem_84_5_W0_addr = W0_addr[25:0];
  assign mem_84_5_W0_clk = W0_clk;
  assign mem_84_5_W0_data = W0_data[47:40];
  assign mem_84_5_W0_en = W0_en & W0_addr_sel == 8'h54;
  assign mem_84_5_W0_mask = W0_mask[5];
  assign mem_84_6_R0_addr = R0_addr[25:0];
  assign mem_84_6_R0_clk = R0_clk;
  assign mem_84_6_R0_en = R0_en & R0_addr_sel == 8'h54;
  assign mem_84_6_W0_addr = W0_addr[25:0];
  assign mem_84_6_W0_clk = W0_clk;
  assign mem_84_6_W0_data = W0_data[55:48];
  assign mem_84_6_W0_en = W0_en & W0_addr_sel == 8'h54;
  assign mem_84_6_W0_mask = W0_mask[6];
  assign mem_84_7_R0_addr = R0_addr[25:0];
  assign mem_84_7_R0_clk = R0_clk;
  assign mem_84_7_R0_en = R0_en & R0_addr_sel == 8'h54;
  assign mem_84_7_W0_addr = W0_addr[25:0];
  assign mem_84_7_W0_clk = W0_clk;
  assign mem_84_7_W0_data = W0_data[63:56];
  assign mem_84_7_W0_en = W0_en & W0_addr_sel == 8'h54;
  assign mem_84_7_W0_mask = W0_mask[7];
  assign mem_85_0_R0_addr = R0_addr[25:0];
  assign mem_85_0_R0_clk = R0_clk;
  assign mem_85_0_R0_en = R0_en & R0_addr_sel == 8'h55;
  assign mem_85_0_W0_addr = W0_addr[25:0];
  assign mem_85_0_W0_clk = W0_clk;
  assign mem_85_0_W0_data = W0_data[7:0];
  assign mem_85_0_W0_en = W0_en & W0_addr_sel == 8'h55;
  assign mem_85_0_W0_mask = W0_mask[0];
  assign mem_85_1_R0_addr = R0_addr[25:0];
  assign mem_85_1_R0_clk = R0_clk;
  assign mem_85_1_R0_en = R0_en & R0_addr_sel == 8'h55;
  assign mem_85_1_W0_addr = W0_addr[25:0];
  assign mem_85_1_W0_clk = W0_clk;
  assign mem_85_1_W0_data = W0_data[15:8];
  assign mem_85_1_W0_en = W0_en & W0_addr_sel == 8'h55;
  assign mem_85_1_W0_mask = W0_mask[1];
  assign mem_85_2_R0_addr = R0_addr[25:0];
  assign mem_85_2_R0_clk = R0_clk;
  assign mem_85_2_R0_en = R0_en & R0_addr_sel == 8'h55;
  assign mem_85_2_W0_addr = W0_addr[25:0];
  assign mem_85_2_W0_clk = W0_clk;
  assign mem_85_2_W0_data = W0_data[23:16];
  assign mem_85_2_W0_en = W0_en & W0_addr_sel == 8'h55;
  assign mem_85_2_W0_mask = W0_mask[2];
  assign mem_85_3_R0_addr = R0_addr[25:0];
  assign mem_85_3_R0_clk = R0_clk;
  assign mem_85_3_R0_en = R0_en & R0_addr_sel == 8'h55;
  assign mem_85_3_W0_addr = W0_addr[25:0];
  assign mem_85_3_W0_clk = W0_clk;
  assign mem_85_3_W0_data = W0_data[31:24];
  assign mem_85_3_W0_en = W0_en & W0_addr_sel == 8'h55;
  assign mem_85_3_W0_mask = W0_mask[3];
  assign mem_85_4_R0_addr = R0_addr[25:0];
  assign mem_85_4_R0_clk = R0_clk;
  assign mem_85_4_R0_en = R0_en & R0_addr_sel == 8'h55;
  assign mem_85_4_W0_addr = W0_addr[25:0];
  assign mem_85_4_W0_clk = W0_clk;
  assign mem_85_4_W0_data = W0_data[39:32];
  assign mem_85_4_W0_en = W0_en & W0_addr_sel == 8'h55;
  assign mem_85_4_W0_mask = W0_mask[4];
  assign mem_85_5_R0_addr = R0_addr[25:0];
  assign mem_85_5_R0_clk = R0_clk;
  assign mem_85_5_R0_en = R0_en & R0_addr_sel == 8'h55;
  assign mem_85_5_W0_addr = W0_addr[25:0];
  assign mem_85_5_W0_clk = W0_clk;
  assign mem_85_5_W0_data = W0_data[47:40];
  assign mem_85_5_W0_en = W0_en & W0_addr_sel == 8'h55;
  assign mem_85_5_W0_mask = W0_mask[5];
  assign mem_85_6_R0_addr = R0_addr[25:0];
  assign mem_85_6_R0_clk = R0_clk;
  assign mem_85_6_R0_en = R0_en & R0_addr_sel == 8'h55;
  assign mem_85_6_W0_addr = W0_addr[25:0];
  assign mem_85_6_W0_clk = W0_clk;
  assign mem_85_6_W0_data = W0_data[55:48];
  assign mem_85_6_W0_en = W0_en & W0_addr_sel == 8'h55;
  assign mem_85_6_W0_mask = W0_mask[6];
  assign mem_85_7_R0_addr = R0_addr[25:0];
  assign mem_85_7_R0_clk = R0_clk;
  assign mem_85_7_R0_en = R0_en & R0_addr_sel == 8'h55;
  assign mem_85_7_W0_addr = W0_addr[25:0];
  assign mem_85_7_W0_clk = W0_clk;
  assign mem_85_7_W0_data = W0_data[63:56];
  assign mem_85_7_W0_en = W0_en & W0_addr_sel == 8'h55;
  assign mem_85_7_W0_mask = W0_mask[7];
  assign mem_86_0_R0_addr = R0_addr[25:0];
  assign mem_86_0_R0_clk = R0_clk;
  assign mem_86_0_R0_en = R0_en & R0_addr_sel == 8'h56;
  assign mem_86_0_W0_addr = W0_addr[25:0];
  assign mem_86_0_W0_clk = W0_clk;
  assign mem_86_0_W0_data = W0_data[7:0];
  assign mem_86_0_W0_en = W0_en & W0_addr_sel == 8'h56;
  assign mem_86_0_W0_mask = W0_mask[0];
  assign mem_86_1_R0_addr = R0_addr[25:0];
  assign mem_86_1_R0_clk = R0_clk;
  assign mem_86_1_R0_en = R0_en & R0_addr_sel == 8'h56;
  assign mem_86_1_W0_addr = W0_addr[25:0];
  assign mem_86_1_W0_clk = W0_clk;
  assign mem_86_1_W0_data = W0_data[15:8];
  assign mem_86_1_W0_en = W0_en & W0_addr_sel == 8'h56;
  assign mem_86_1_W0_mask = W0_mask[1];
  assign mem_86_2_R0_addr = R0_addr[25:0];
  assign mem_86_2_R0_clk = R0_clk;
  assign mem_86_2_R0_en = R0_en & R0_addr_sel == 8'h56;
  assign mem_86_2_W0_addr = W0_addr[25:0];
  assign mem_86_2_W0_clk = W0_clk;
  assign mem_86_2_W0_data = W0_data[23:16];
  assign mem_86_2_W0_en = W0_en & W0_addr_sel == 8'h56;
  assign mem_86_2_W0_mask = W0_mask[2];
  assign mem_86_3_R0_addr = R0_addr[25:0];
  assign mem_86_3_R0_clk = R0_clk;
  assign mem_86_3_R0_en = R0_en & R0_addr_sel == 8'h56;
  assign mem_86_3_W0_addr = W0_addr[25:0];
  assign mem_86_3_W0_clk = W0_clk;
  assign mem_86_3_W0_data = W0_data[31:24];
  assign mem_86_3_W0_en = W0_en & W0_addr_sel == 8'h56;
  assign mem_86_3_W0_mask = W0_mask[3];
  assign mem_86_4_R0_addr = R0_addr[25:0];
  assign mem_86_4_R0_clk = R0_clk;
  assign mem_86_4_R0_en = R0_en & R0_addr_sel == 8'h56;
  assign mem_86_4_W0_addr = W0_addr[25:0];
  assign mem_86_4_W0_clk = W0_clk;
  assign mem_86_4_W0_data = W0_data[39:32];
  assign mem_86_4_W0_en = W0_en & W0_addr_sel == 8'h56;
  assign mem_86_4_W0_mask = W0_mask[4];
  assign mem_86_5_R0_addr = R0_addr[25:0];
  assign mem_86_5_R0_clk = R0_clk;
  assign mem_86_5_R0_en = R0_en & R0_addr_sel == 8'h56;
  assign mem_86_5_W0_addr = W0_addr[25:0];
  assign mem_86_5_W0_clk = W0_clk;
  assign mem_86_5_W0_data = W0_data[47:40];
  assign mem_86_5_W0_en = W0_en & W0_addr_sel == 8'h56;
  assign mem_86_5_W0_mask = W0_mask[5];
  assign mem_86_6_R0_addr = R0_addr[25:0];
  assign mem_86_6_R0_clk = R0_clk;
  assign mem_86_6_R0_en = R0_en & R0_addr_sel == 8'h56;
  assign mem_86_6_W0_addr = W0_addr[25:0];
  assign mem_86_6_W0_clk = W0_clk;
  assign mem_86_6_W0_data = W0_data[55:48];
  assign mem_86_6_W0_en = W0_en & W0_addr_sel == 8'h56;
  assign mem_86_6_W0_mask = W0_mask[6];
  assign mem_86_7_R0_addr = R0_addr[25:0];
  assign mem_86_7_R0_clk = R0_clk;
  assign mem_86_7_R0_en = R0_en & R0_addr_sel == 8'h56;
  assign mem_86_7_W0_addr = W0_addr[25:0];
  assign mem_86_7_W0_clk = W0_clk;
  assign mem_86_7_W0_data = W0_data[63:56];
  assign mem_86_7_W0_en = W0_en & W0_addr_sel == 8'h56;
  assign mem_86_7_W0_mask = W0_mask[7];
  assign mem_87_0_R0_addr = R0_addr[25:0];
  assign mem_87_0_R0_clk = R0_clk;
  assign mem_87_0_R0_en = R0_en & R0_addr_sel == 8'h57;
  assign mem_87_0_W0_addr = W0_addr[25:0];
  assign mem_87_0_W0_clk = W0_clk;
  assign mem_87_0_W0_data = W0_data[7:0];
  assign mem_87_0_W0_en = W0_en & W0_addr_sel == 8'h57;
  assign mem_87_0_W0_mask = W0_mask[0];
  assign mem_87_1_R0_addr = R0_addr[25:0];
  assign mem_87_1_R0_clk = R0_clk;
  assign mem_87_1_R0_en = R0_en & R0_addr_sel == 8'h57;
  assign mem_87_1_W0_addr = W0_addr[25:0];
  assign mem_87_1_W0_clk = W0_clk;
  assign mem_87_1_W0_data = W0_data[15:8];
  assign mem_87_1_W0_en = W0_en & W0_addr_sel == 8'h57;
  assign mem_87_1_W0_mask = W0_mask[1];
  assign mem_87_2_R0_addr = R0_addr[25:0];
  assign mem_87_2_R0_clk = R0_clk;
  assign mem_87_2_R0_en = R0_en & R0_addr_sel == 8'h57;
  assign mem_87_2_W0_addr = W0_addr[25:0];
  assign mem_87_2_W0_clk = W0_clk;
  assign mem_87_2_W0_data = W0_data[23:16];
  assign mem_87_2_W0_en = W0_en & W0_addr_sel == 8'h57;
  assign mem_87_2_W0_mask = W0_mask[2];
  assign mem_87_3_R0_addr = R0_addr[25:0];
  assign mem_87_3_R0_clk = R0_clk;
  assign mem_87_3_R0_en = R0_en & R0_addr_sel == 8'h57;
  assign mem_87_3_W0_addr = W0_addr[25:0];
  assign mem_87_3_W0_clk = W0_clk;
  assign mem_87_3_W0_data = W0_data[31:24];
  assign mem_87_3_W0_en = W0_en & W0_addr_sel == 8'h57;
  assign mem_87_3_W0_mask = W0_mask[3];
  assign mem_87_4_R0_addr = R0_addr[25:0];
  assign mem_87_4_R0_clk = R0_clk;
  assign mem_87_4_R0_en = R0_en & R0_addr_sel == 8'h57;
  assign mem_87_4_W0_addr = W0_addr[25:0];
  assign mem_87_4_W0_clk = W0_clk;
  assign mem_87_4_W0_data = W0_data[39:32];
  assign mem_87_4_W0_en = W0_en & W0_addr_sel == 8'h57;
  assign mem_87_4_W0_mask = W0_mask[4];
  assign mem_87_5_R0_addr = R0_addr[25:0];
  assign mem_87_5_R0_clk = R0_clk;
  assign mem_87_5_R0_en = R0_en & R0_addr_sel == 8'h57;
  assign mem_87_5_W0_addr = W0_addr[25:0];
  assign mem_87_5_W0_clk = W0_clk;
  assign mem_87_5_W0_data = W0_data[47:40];
  assign mem_87_5_W0_en = W0_en & W0_addr_sel == 8'h57;
  assign mem_87_5_W0_mask = W0_mask[5];
  assign mem_87_6_R0_addr = R0_addr[25:0];
  assign mem_87_6_R0_clk = R0_clk;
  assign mem_87_6_R0_en = R0_en & R0_addr_sel == 8'h57;
  assign mem_87_6_W0_addr = W0_addr[25:0];
  assign mem_87_6_W0_clk = W0_clk;
  assign mem_87_6_W0_data = W0_data[55:48];
  assign mem_87_6_W0_en = W0_en & W0_addr_sel == 8'h57;
  assign mem_87_6_W0_mask = W0_mask[6];
  assign mem_87_7_R0_addr = R0_addr[25:0];
  assign mem_87_7_R0_clk = R0_clk;
  assign mem_87_7_R0_en = R0_en & R0_addr_sel == 8'h57;
  assign mem_87_7_W0_addr = W0_addr[25:0];
  assign mem_87_7_W0_clk = W0_clk;
  assign mem_87_7_W0_data = W0_data[63:56];
  assign mem_87_7_W0_en = W0_en & W0_addr_sel == 8'h57;
  assign mem_87_7_W0_mask = W0_mask[7];
  assign mem_88_0_R0_addr = R0_addr[25:0];
  assign mem_88_0_R0_clk = R0_clk;
  assign mem_88_0_R0_en = R0_en & R0_addr_sel == 8'h58;
  assign mem_88_0_W0_addr = W0_addr[25:0];
  assign mem_88_0_W0_clk = W0_clk;
  assign mem_88_0_W0_data = W0_data[7:0];
  assign mem_88_0_W0_en = W0_en & W0_addr_sel == 8'h58;
  assign mem_88_0_W0_mask = W0_mask[0];
  assign mem_88_1_R0_addr = R0_addr[25:0];
  assign mem_88_1_R0_clk = R0_clk;
  assign mem_88_1_R0_en = R0_en & R0_addr_sel == 8'h58;
  assign mem_88_1_W0_addr = W0_addr[25:0];
  assign mem_88_1_W0_clk = W0_clk;
  assign mem_88_1_W0_data = W0_data[15:8];
  assign mem_88_1_W0_en = W0_en & W0_addr_sel == 8'h58;
  assign mem_88_1_W0_mask = W0_mask[1];
  assign mem_88_2_R0_addr = R0_addr[25:0];
  assign mem_88_2_R0_clk = R0_clk;
  assign mem_88_2_R0_en = R0_en & R0_addr_sel == 8'h58;
  assign mem_88_2_W0_addr = W0_addr[25:0];
  assign mem_88_2_W0_clk = W0_clk;
  assign mem_88_2_W0_data = W0_data[23:16];
  assign mem_88_2_W0_en = W0_en & W0_addr_sel == 8'h58;
  assign mem_88_2_W0_mask = W0_mask[2];
  assign mem_88_3_R0_addr = R0_addr[25:0];
  assign mem_88_3_R0_clk = R0_clk;
  assign mem_88_3_R0_en = R0_en & R0_addr_sel == 8'h58;
  assign mem_88_3_W0_addr = W0_addr[25:0];
  assign mem_88_3_W0_clk = W0_clk;
  assign mem_88_3_W0_data = W0_data[31:24];
  assign mem_88_3_W0_en = W0_en & W0_addr_sel == 8'h58;
  assign mem_88_3_W0_mask = W0_mask[3];
  assign mem_88_4_R0_addr = R0_addr[25:0];
  assign mem_88_4_R0_clk = R0_clk;
  assign mem_88_4_R0_en = R0_en & R0_addr_sel == 8'h58;
  assign mem_88_4_W0_addr = W0_addr[25:0];
  assign mem_88_4_W0_clk = W0_clk;
  assign mem_88_4_W0_data = W0_data[39:32];
  assign mem_88_4_W0_en = W0_en & W0_addr_sel == 8'h58;
  assign mem_88_4_W0_mask = W0_mask[4];
  assign mem_88_5_R0_addr = R0_addr[25:0];
  assign mem_88_5_R0_clk = R0_clk;
  assign mem_88_5_R0_en = R0_en & R0_addr_sel == 8'h58;
  assign mem_88_5_W0_addr = W0_addr[25:0];
  assign mem_88_5_W0_clk = W0_clk;
  assign mem_88_5_W0_data = W0_data[47:40];
  assign mem_88_5_W0_en = W0_en & W0_addr_sel == 8'h58;
  assign mem_88_5_W0_mask = W0_mask[5];
  assign mem_88_6_R0_addr = R0_addr[25:0];
  assign mem_88_6_R0_clk = R0_clk;
  assign mem_88_6_R0_en = R0_en & R0_addr_sel == 8'h58;
  assign mem_88_6_W0_addr = W0_addr[25:0];
  assign mem_88_6_W0_clk = W0_clk;
  assign mem_88_6_W0_data = W0_data[55:48];
  assign mem_88_6_W0_en = W0_en & W0_addr_sel == 8'h58;
  assign mem_88_6_W0_mask = W0_mask[6];
  assign mem_88_7_R0_addr = R0_addr[25:0];
  assign mem_88_7_R0_clk = R0_clk;
  assign mem_88_7_R0_en = R0_en & R0_addr_sel == 8'h58;
  assign mem_88_7_W0_addr = W0_addr[25:0];
  assign mem_88_7_W0_clk = W0_clk;
  assign mem_88_7_W0_data = W0_data[63:56];
  assign mem_88_7_W0_en = W0_en & W0_addr_sel == 8'h58;
  assign mem_88_7_W0_mask = W0_mask[7];
  assign mem_89_0_R0_addr = R0_addr[25:0];
  assign mem_89_0_R0_clk = R0_clk;
  assign mem_89_0_R0_en = R0_en & R0_addr_sel == 8'h59;
  assign mem_89_0_W0_addr = W0_addr[25:0];
  assign mem_89_0_W0_clk = W0_clk;
  assign mem_89_0_W0_data = W0_data[7:0];
  assign mem_89_0_W0_en = W0_en & W0_addr_sel == 8'h59;
  assign mem_89_0_W0_mask = W0_mask[0];
  assign mem_89_1_R0_addr = R0_addr[25:0];
  assign mem_89_1_R0_clk = R0_clk;
  assign mem_89_1_R0_en = R0_en & R0_addr_sel == 8'h59;
  assign mem_89_1_W0_addr = W0_addr[25:0];
  assign mem_89_1_W0_clk = W0_clk;
  assign mem_89_1_W0_data = W0_data[15:8];
  assign mem_89_1_W0_en = W0_en & W0_addr_sel == 8'h59;
  assign mem_89_1_W0_mask = W0_mask[1];
  assign mem_89_2_R0_addr = R0_addr[25:0];
  assign mem_89_2_R0_clk = R0_clk;
  assign mem_89_2_R0_en = R0_en & R0_addr_sel == 8'h59;
  assign mem_89_2_W0_addr = W0_addr[25:0];
  assign mem_89_2_W0_clk = W0_clk;
  assign mem_89_2_W0_data = W0_data[23:16];
  assign mem_89_2_W0_en = W0_en & W0_addr_sel == 8'h59;
  assign mem_89_2_W0_mask = W0_mask[2];
  assign mem_89_3_R0_addr = R0_addr[25:0];
  assign mem_89_3_R0_clk = R0_clk;
  assign mem_89_3_R0_en = R0_en & R0_addr_sel == 8'h59;
  assign mem_89_3_W0_addr = W0_addr[25:0];
  assign mem_89_3_W0_clk = W0_clk;
  assign mem_89_3_W0_data = W0_data[31:24];
  assign mem_89_3_W0_en = W0_en & W0_addr_sel == 8'h59;
  assign mem_89_3_W0_mask = W0_mask[3];
  assign mem_89_4_R0_addr = R0_addr[25:0];
  assign mem_89_4_R0_clk = R0_clk;
  assign mem_89_4_R0_en = R0_en & R0_addr_sel == 8'h59;
  assign mem_89_4_W0_addr = W0_addr[25:0];
  assign mem_89_4_W0_clk = W0_clk;
  assign mem_89_4_W0_data = W0_data[39:32];
  assign mem_89_4_W0_en = W0_en & W0_addr_sel == 8'h59;
  assign mem_89_4_W0_mask = W0_mask[4];
  assign mem_89_5_R0_addr = R0_addr[25:0];
  assign mem_89_5_R0_clk = R0_clk;
  assign mem_89_5_R0_en = R0_en & R0_addr_sel == 8'h59;
  assign mem_89_5_W0_addr = W0_addr[25:0];
  assign mem_89_5_W0_clk = W0_clk;
  assign mem_89_5_W0_data = W0_data[47:40];
  assign mem_89_5_W0_en = W0_en & W0_addr_sel == 8'h59;
  assign mem_89_5_W0_mask = W0_mask[5];
  assign mem_89_6_R0_addr = R0_addr[25:0];
  assign mem_89_6_R0_clk = R0_clk;
  assign mem_89_6_R0_en = R0_en & R0_addr_sel == 8'h59;
  assign mem_89_6_W0_addr = W0_addr[25:0];
  assign mem_89_6_W0_clk = W0_clk;
  assign mem_89_6_W0_data = W0_data[55:48];
  assign mem_89_6_W0_en = W0_en & W0_addr_sel == 8'h59;
  assign mem_89_6_W0_mask = W0_mask[6];
  assign mem_89_7_R0_addr = R0_addr[25:0];
  assign mem_89_7_R0_clk = R0_clk;
  assign mem_89_7_R0_en = R0_en & R0_addr_sel == 8'h59;
  assign mem_89_7_W0_addr = W0_addr[25:0];
  assign mem_89_7_W0_clk = W0_clk;
  assign mem_89_7_W0_data = W0_data[63:56];
  assign mem_89_7_W0_en = W0_en & W0_addr_sel == 8'h59;
  assign mem_89_7_W0_mask = W0_mask[7];
  assign mem_90_0_R0_addr = R0_addr[25:0];
  assign mem_90_0_R0_clk = R0_clk;
  assign mem_90_0_R0_en = R0_en & R0_addr_sel == 8'h5a;
  assign mem_90_0_W0_addr = W0_addr[25:0];
  assign mem_90_0_W0_clk = W0_clk;
  assign mem_90_0_W0_data = W0_data[7:0];
  assign mem_90_0_W0_en = W0_en & W0_addr_sel == 8'h5a;
  assign mem_90_0_W0_mask = W0_mask[0];
  assign mem_90_1_R0_addr = R0_addr[25:0];
  assign mem_90_1_R0_clk = R0_clk;
  assign mem_90_1_R0_en = R0_en & R0_addr_sel == 8'h5a;
  assign mem_90_1_W0_addr = W0_addr[25:0];
  assign mem_90_1_W0_clk = W0_clk;
  assign mem_90_1_W0_data = W0_data[15:8];
  assign mem_90_1_W0_en = W0_en & W0_addr_sel == 8'h5a;
  assign mem_90_1_W0_mask = W0_mask[1];
  assign mem_90_2_R0_addr = R0_addr[25:0];
  assign mem_90_2_R0_clk = R0_clk;
  assign mem_90_2_R0_en = R0_en & R0_addr_sel == 8'h5a;
  assign mem_90_2_W0_addr = W0_addr[25:0];
  assign mem_90_2_W0_clk = W0_clk;
  assign mem_90_2_W0_data = W0_data[23:16];
  assign mem_90_2_W0_en = W0_en & W0_addr_sel == 8'h5a;
  assign mem_90_2_W0_mask = W0_mask[2];
  assign mem_90_3_R0_addr = R0_addr[25:0];
  assign mem_90_3_R0_clk = R0_clk;
  assign mem_90_3_R0_en = R0_en & R0_addr_sel == 8'h5a;
  assign mem_90_3_W0_addr = W0_addr[25:0];
  assign mem_90_3_W0_clk = W0_clk;
  assign mem_90_3_W0_data = W0_data[31:24];
  assign mem_90_3_W0_en = W0_en & W0_addr_sel == 8'h5a;
  assign mem_90_3_W0_mask = W0_mask[3];
  assign mem_90_4_R0_addr = R0_addr[25:0];
  assign mem_90_4_R0_clk = R0_clk;
  assign mem_90_4_R0_en = R0_en & R0_addr_sel == 8'h5a;
  assign mem_90_4_W0_addr = W0_addr[25:0];
  assign mem_90_4_W0_clk = W0_clk;
  assign mem_90_4_W0_data = W0_data[39:32];
  assign mem_90_4_W0_en = W0_en & W0_addr_sel == 8'h5a;
  assign mem_90_4_W0_mask = W0_mask[4];
  assign mem_90_5_R0_addr = R0_addr[25:0];
  assign mem_90_5_R0_clk = R0_clk;
  assign mem_90_5_R0_en = R0_en & R0_addr_sel == 8'h5a;
  assign mem_90_5_W0_addr = W0_addr[25:0];
  assign mem_90_5_W0_clk = W0_clk;
  assign mem_90_5_W0_data = W0_data[47:40];
  assign mem_90_5_W0_en = W0_en & W0_addr_sel == 8'h5a;
  assign mem_90_5_W0_mask = W0_mask[5];
  assign mem_90_6_R0_addr = R0_addr[25:0];
  assign mem_90_6_R0_clk = R0_clk;
  assign mem_90_6_R0_en = R0_en & R0_addr_sel == 8'h5a;
  assign mem_90_6_W0_addr = W0_addr[25:0];
  assign mem_90_6_W0_clk = W0_clk;
  assign mem_90_6_W0_data = W0_data[55:48];
  assign mem_90_6_W0_en = W0_en & W0_addr_sel == 8'h5a;
  assign mem_90_6_W0_mask = W0_mask[6];
  assign mem_90_7_R0_addr = R0_addr[25:0];
  assign mem_90_7_R0_clk = R0_clk;
  assign mem_90_7_R0_en = R0_en & R0_addr_sel == 8'h5a;
  assign mem_90_7_W0_addr = W0_addr[25:0];
  assign mem_90_7_W0_clk = W0_clk;
  assign mem_90_7_W0_data = W0_data[63:56];
  assign mem_90_7_W0_en = W0_en & W0_addr_sel == 8'h5a;
  assign mem_90_7_W0_mask = W0_mask[7];
  assign mem_91_0_R0_addr = R0_addr[25:0];
  assign mem_91_0_R0_clk = R0_clk;
  assign mem_91_0_R0_en = R0_en & R0_addr_sel == 8'h5b;
  assign mem_91_0_W0_addr = W0_addr[25:0];
  assign mem_91_0_W0_clk = W0_clk;
  assign mem_91_0_W0_data = W0_data[7:0];
  assign mem_91_0_W0_en = W0_en & W0_addr_sel == 8'h5b;
  assign mem_91_0_W0_mask = W0_mask[0];
  assign mem_91_1_R0_addr = R0_addr[25:0];
  assign mem_91_1_R0_clk = R0_clk;
  assign mem_91_1_R0_en = R0_en & R0_addr_sel == 8'h5b;
  assign mem_91_1_W0_addr = W0_addr[25:0];
  assign mem_91_1_W0_clk = W0_clk;
  assign mem_91_1_W0_data = W0_data[15:8];
  assign mem_91_1_W0_en = W0_en & W0_addr_sel == 8'h5b;
  assign mem_91_1_W0_mask = W0_mask[1];
  assign mem_91_2_R0_addr = R0_addr[25:0];
  assign mem_91_2_R0_clk = R0_clk;
  assign mem_91_2_R0_en = R0_en & R0_addr_sel == 8'h5b;
  assign mem_91_2_W0_addr = W0_addr[25:0];
  assign mem_91_2_W0_clk = W0_clk;
  assign mem_91_2_W0_data = W0_data[23:16];
  assign mem_91_2_W0_en = W0_en & W0_addr_sel == 8'h5b;
  assign mem_91_2_W0_mask = W0_mask[2];
  assign mem_91_3_R0_addr = R0_addr[25:0];
  assign mem_91_3_R0_clk = R0_clk;
  assign mem_91_3_R0_en = R0_en & R0_addr_sel == 8'h5b;
  assign mem_91_3_W0_addr = W0_addr[25:0];
  assign mem_91_3_W0_clk = W0_clk;
  assign mem_91_3_W0_data = W0_data[31:24];
  assign mem_91_3_W0_en = W0_en & W0_addr_sel == 8'h5b;
  assign mem_91_3_W0_mask = W0_mask[3];
  assign mem_91_4_R0_addr = R0_addr[25:0];
  assign mem_91_4_R0_clk = R0_clk;
  assign mem_91_4_R0_en = R0_en & R0_addr_sel == 8'h5b;
  assign mem_91_4_W0_addr = W0_addr[25:0];
  assign mem_91_4_W0_clk = W0_clk;
  assign mem_91_4_W0_data = W0_data[39:32];
  assign mem_91_4_W0_en = W0_en & W0_addr_sel == 8'h5b;
  assign mem_91_4_W0_mask = W0_mask[4];
  assign mem_91_5_R0_addr = R0_addr[25:0];
  assign mem_91_5_R0_clk = R0_clk;
  assign mem_91_5_R0_en = R0_en & R0_addr_sel == 8'h5b;
  assign mem_91_5_W0_addr = W0_addr[25:0];
  assign mem_91_5_W0_clk = W0_clk;
  assign mem_91_5_W0_data = W0_data[47:40];
  assign mem_91_5_W0_en = W0_en & W0_addr_sel == 8'h5b;
  assign mem_91_5_W0_mask = W0_mask[5];
  assign mem_91_6_R0_addr = R0_addr[25:0];
  assign mem_91_6_R0_clk = R0_clk;
  assign mem_91_6_R0_en = R0_en & R0_addr_sel == 8'h5b;
  assign mem_91_6_W0_addr = W0_addr[25:0];
  assign mem_91_6_W0_clk = W0_clk;
  assign mem_91_6_W0_data = W0_data[55:48];
  assign mem_91_6_W0_en = W0_en & W0_addr_sel == 8'h5b;
  assign mem_91_6_W0_mask = W0_mask[6];
  assign mem_91_7_R0_addr = R0_addr[25:0];
  assign mem_91_7_R0_clk = R0_clk;
  assign mem_91_7_R0_en = R0_en & R0_addr_sel == 8'h5b;
  assign mem_91_7_W0_addr = W0_addr[25:0];
  assign mem_91_7_W0_clk = W0_clk;
  assign mem_91_7_W0_data = W0_data[63:56];
  assign mem_91_7_W0_en = W0_en & W0_addr_sel == 8'h5b;
  assign mem_91_7_W0_mask = W0_mask[7];
  assign mem_92_0_R0_addr = R0_addr[25:0];
  assign mem_92_0_R0_clk = R0_clk;
  assign mem_92_0_R0_en = R0_en & R0_addr_sel == 8'h5c;
  assign mem_92_0_W0_addr = W0_addr[25:0];
  assign mem_92_0_W0_clk = W0_clk;
  assign mem_92_0_W0_data = W0_data[7:0];
  assign mem_92_0_W0_en = W0_en & W0_addr_sel == 8'h5c;
  assign mem_92_0_W0_mask = W0_mask[0];
  assign mem_92_1_R0_addr = R0_addr[25:0];
  assign mem_92_1_R0_clk = R0_clk;
  assign mem_92_1_R0_en = R0_en & R0_addr_sel == 8'h5c;
  assign mem_92_1_W0_addr = W0_addr[25:0];
  assign mem_92_1_W0_clk = W0_clk;
  assign mem_92_1_W0_data = W0_data[15:8];
  assign mem_92_1_W0_en = W0_en & W0_addr_sel == 8'h5c;
  assign mem_92_1_W0_mask = W0_mask[1];
  assign mem_92_2_R0_addr = R0_addr[25:0];
  assign mem_92_2_R0_clk = R0_clk;
  assign mem_92_2_R0_en = R0_en & R0_addr_sel == 8'h5c;
  assign mem_92_2_W0_addr = W0_addr[25:0];
  assign mem_92_2_W0_clk = W0_clk;
  assign mem_92_2_W0_data = W0_data[23:16];
  assign mem_92_2_W0_en = W0_en & W0_addr_sel == 8'h5c;
  assign mem_92_2_W0_mask = W0_mask[2];
  assign mem_92_3_R0_addr = R0_addr[25:0];
  assign mem_92_3_R0_clk = R0_clk;
  assign mem_92_3_R0_en = R0_en & R0_addr_sel == 8'h5c;
  assign mem_92_3_W0_addr = W0_addr[25:0];
  assign mem_92_3_W0_clk = W0_clk;
  assign mem_92_3_W0_data = W0_data[31:24];
  assign mem_92_3_W0_en = W0_en & W0_addr_sel == 8'h5c;
  assign mem_92_3_W0_mask = W0_mask[3];
  assign mem_92_4_R0_addr = R0_addr[25:0];
  assign mem_92_4_R0_clk = R0_clk;
  assign mem_92_4_R0_en = R0_en & R0_addr_sel == 8'h5c;
  assign mem_92_4_W0_addr = W0_addr[25:0];
  assign mem_92_4_W0_clk = W0_clk;
  assign mem_92_4_W0_data = W0_data[39:32];
  assign mem_92_4_W0_en = W0_en & W0_addr_sel == 8'h5c;
  assign mem_92_4_W0_mask = W0_mask[4];
  assign mem_92_5_R0_addr = R0_addr[25:0];
  assign mem_92_5_R0_clk = R0_clk;
  assign mem_92_5_R0_en = R0_en & R0_addr_sel == 8'h5c;
  assign mem_92_5_W0_addr = W0_addr[25:0];
  assign mem_92_5_W0_clk = W0_clk;
  assign mem_92_5_W0_data = W0_data[47:40];
  assign mem_92_5_W0_en = W0_en & W0_addr_sel == 8'h5c;
  assign mem_92_5_W0_mask = W0_mask[5];
  assign mem_92_6_R0_addr = R0_addr[25:0];
  assign mem_92_6_R0_clk = R0_clk;
  assign mem_92_6_R0_en = R0_en & R0_addr_sel == 8'h5c;
  assign mem_92_6_W0_addr = W0_addr[25:0];
  assign mem_92_6_W0_clk = W0_clk;
  assign mem_92_6_W0_data = W0_data[55:48];
  assign mem_92_6_W0_en = W0_en & W0_addr_sel == 8'h5c;
  assign mem_92_6_W0_mask = W0_mask[6];
  assign mem_92_7_R0_addr = R0_addr[25:0];
  assign mem_92_7_R0_clk = R0_clk;
  assign mem_92_7_R0_en = R0_en & R0_addr_sel == 8'h5c;
  assign mem_92_7_W0_addr = W0_addr[25:0];
  assign mem_92_7_W0_clk = W0_clk;
  assign mem_92_7_W0_data = W0_data[63:56];
  assign mem_92_7_W0_en = W0_en & W0_addr_sel == 8'h5c;
  assign mem_92_7_W0_mask = W0_mask[7];
  assign mem_93_0_R0_addr = R0_addr[25:0];
  assign mem_93_0_R0_clk = R0_clk;
  assign mem_93_0_R0_en = R0_en & R0_addr_sel == 8'h5d;
  assign mem_93_0_W0_addr = W0_addr[25:0];
  assign mem_93_0_W0_clk = W0_clk;
  assign mem_93_0_W0_data = W0_data[7:0];
  assign mem_93_0_W0_en = W0_en & W0_addr_sel == 8'h5d;
  assign mem_93_0_W0_mask = W0_mask[0];
  assign mem_93_1_R0_addr = R0_addr[25:0];
  assign mem_93_1_R0_clk = R0_clk;
  assign mem_93_1_R0_en = R0_en & R0_addr_sel == 8'h5d;
  assign mem_93_1_W0_addr = W0_addr[25:0];
  assign mem_93_1_W0_clk = W0_clk;
  assign mem_93_1_W0_data = W0_data[15:8];
  assign mem_93_1_W0_en = W0_en & W0_addr_sel == 8'h5d;
  assign mem_93_1_W0_mask = W0_mask[1];
  assign mem_93_2_R0_addr = R0_addr[25:0];
  assign mem_93_2_R0_clk = R0_clk;
  assign mem_93_2_R0_en = R0_en & R0_addr_sel == 8'h5d;
  assign mem_93_2_W0_addr = W0_addr[25:0];
  assign mem_93_2_W0_clk = W0_clk;
  assign mem_93_2_W0_data = W0_data[23:16];
  assign mem_93_2_W0_en = W0_en & W0_addr_sel == 8'h5d;
  assign mem_93_2_W0_mask = W0_mask[2];
  assign mem_93_3_R0_addr = R0_addr[25:0];
  assign mem_93_3_R0_clk = R0_clk;
  assign mem_93_3_R0_en = R0_en & R0_addr_sel == 8'h5d;
  assign mem_93_3_W0_addr = W0_addr[25:0];
  assign mem_93_3_W0_clk = W0_clk;
  assign mem_93_3_W0_data = W0_data[31:24];
  assign mem_93_3_W0_en = W0_en & W0_addr_sel == 8'h5d;
  assign mem_93_3_W0_mask = W0_mask[3];
  assign mem_93_4_R0_addr = R0_addr[25:0];
  assign mem_93_4_R0_clk = R0_clk;
  assign mem_93_4_R0_en = R0_en & R0_addr_sel == 8'h5d;
  assign mem_93_4_W0_addr = W0_addr[25:0];
  assign mem_93_4_W0_clk = W0_clk;
  assign mem_93_4_W0_data = W0_data[39:32];
  assign mem_93_4_W0_en = W0_en & W0_addr_sel == 8'h5d;
  assign mem_93_4_W0_mask = W0_mask[4];
  assign mem_93_5_R0_addr = R0_addr[25:0];
  assign mem_93_5_R0_clk = R0_clk;
  assign mem_93_5_R0_en = R0_en & R0_addr_sel == 8'h5d;
  assign mem_93_5_W0_addr = W0_addr[25:0];
  assign mem_93_5_W0_clk = W0_clk;
  assign mem_93_5_W0_data = W0_data[47:40];
  assign mem_93_5_W0_en = W0_en & W0_addr_sel == 8'h5d;
  assign mem_93_5_W0_mask = W0_mask[5];
  assign mem_93_6_R0_addr = R0_addr[25:0];
  assign mem_93_6_R0_clk = R0_clk;
  assign mem_93_6_R0_en = R0_en & R0_addr_sel == 8'h5d;
  assign mem_93_6_W0_addr = W0_addr[25:0];
  assign mem_93_6_W0_clk = W0_clk;
  assign mem_93_6_W0_data = W0_data[55:48];
  assign mem_93_6_W0_en = W0_en & W0_addr_sel == 8'h5d;
  assign mem_93_6_W0_mask = W0_mask[6];
  assign mem_93_7_R0_addr = R0_addr[25:0];
  assign mem_93_7_R0_clk = R0_clk;
  assign mem_93_7_R0_en = R0_en & R0_addr_sel == 8'h5d;
  assign mem_93_7_W0_addr = W0_addr[25:0];
  assign mem_93_7_W0_clk = W0_clk;
  assign mem_93_7_W0_data = W0_data[63:56];
  assign mem_93_7_W0_en = W0_en & W0_addr_sel == 8'h5d;
  assign mem_93_7_W0_mask = W0_mask[7];
  assign mem_94_0_R0_addr = R0_addr[25:0];
  assign mem_94_0_R0_clk = R0_clk;
  assign mem_94_0_R0_en = R0_en & R0_addr_sel == 8'h5e;
  assign mem_94_0_W0_addr = W0_addr[25:0];
  assign mem_94_0_W0_clk = W0_clk;
  assign mem_94_0_W0_data = W0_data[7:0];
  assign mem_94_0_W0_en = W0_en & W0_addr_sel == 8'h5e;
  assign mem_94_0_W0_mask = W0_mask[0];
  assign mem_94_1_R0_addr = R0_addr[25:0];
  assign mem_94_1_R0_clk = R0_clk;
  assign mem_94_1_R0_en = R0_en & R0_addr_sel == 8'h5e;
  assign mem_94_1_W0_addr = W0_addr[25:0];
  assign mem_94_1_W0_clk = W0_clk;
  assign mem_94_1_W0_data = W0_data[15:8];
  assign mem_94_1_W0_en = W0_en & W0_addr_sel == 8'h5e;
  assign mem_94_1_W0_mask = W0_mask[1];
  assign mem_94_2_R0_addr = R0_addr[25:0];
  assign mem_94_2_R0_clk = R0_clk;
  assign mem_94_2_R0_en = R0_en & R0_addr_sel == 8'h5e;
  assign mem_94_2_W0_addr = W0_addr[25:0];
  assign mem_94_2_W0_clk = W0_clk;
  assign mem_94_2_W0_data = W0_data[23:16];
  assign mem_94_2_W0_en = W0_en & W0_addr_sel == 8'h5e;
  assign mem_94_2_W0_mask = W0_mask[2];
  assign mem_94_3_R0_addr = R0_addr[25:0];
  assign mem_94_3_R0_clk = R0_clk;
  assign mem_94_3_R0_en = R0_en & R0_addr_sel == 8'h5e;
  assign mem_94_3_W0_addr = W0_addr[25:0];
  assign mem_94_3_W0_clk = W0_clk;
  assign mem_94_3_W0_data = W0_data[31:24];
  assign mem_94_3_W0_en = W0_en & W0_addr_sel == 8'h5e;
  assign mem_94_3_W0_mask = W0_mask[3];
  assign mem_94_4_R0_addr = R0_addr[25:0];
  assign mem_94_4_R0_clk = R0_clk;
  assign mem_94_4_R0_en = R0_en & R0_addr_sel == 8'h5e;
  assign mem_94_4_W0_addr = W0_addr[25:0];
  assign mem_94_4_W0_clk = W0_clk;
  assign mem_94_4_W0_data = W0_data[39:32];
  assign mem_94_4_W0_en = W0_en & W0_addr_sel == 8'h5e;
  assign mem_94_4_W0_mask = W0_mask[4];
  assign mem_94_5_R0_addr = R0_addr[25:0];
  assign mem_94_5_R0_clk = R0_clk;
  assign mem_94_5_R0_en = R0_en & R0_addr_sel == 8'h5e;
  assign mem_94_5_W0_addr = W0_addr[25:0];
  assign mem_94_5_W0_clk = W0_clk;
  assign mem_94_5_W0_data = W0_data[47:40];
  assign mem_94_5_W0_en = W0_en & W0_addr_sel == 8'h5e;
  assign mem_94_5_W0_mask = W0_mask[5];
  assign mem_94_6_R0_addr = R0_addr[25:0];
  assign mem_94_6_R0_clk = R0_clk;
  assign mem_94_6_R0_en = R0_en & R0_addr_sel == 8'h5e;
  assign mem_94_6_W0_addr = W0_addr[25:0];
  assign mem_94_6_W0_clk = W0_clk;
  assign mem_94_6_W0_data = W0_data[55:48];
  assign mem_94_6_W0_en = W0_en & W0_addr_sel == 8'h5e;
  assign mem_94_6_W0_mask = W0_mask[6];
  assign mem_94_7_R0_addr = R0_addr[25:0];
  assign mem_94_7_R0_clk = R0_clk;
  assign mem_94_7_R0_en = R0_en & R0_addr_sel == 8'h5e;
  assign mem_94_7_W0_addr = W0_addr[25:0];
  assign mem_94_7_W0_clk = W0_clk;
  assign mem_94_7_W0_data = W0_data[63:56];
  assign mem_94_7_W0_en = W0_en & W0_addr_sel == 8'h5e;
  assign mem_94_7_W0_mask = W0_mask[7];
  assign mem_95_0_R0_addr = R0_addr[25:0];
  assign mem_95_0_R0_clk = R0_clk;
  assign mem_95_0_R0_en = R0_en & R0_addr_sel == 8'h5f;
  assign mem_95_0_W0_addr = W0_addr[25:0];
  assign mem_95_0_W0_clk = W0_clk;
  assign mem_95_0_W0_data = W0_data[7:0];
  assign mem_95_0_W0_en = W0_en & W0_addr_sel == 8'h5f;
  assign mem_95_0_W0_mask = W0_mask[0];
  assign mem_95_1_R0_addr = R0_addr[25:0];
  assign mem_95_1_R0_clk = R0_clk;
  assign mem_95_1_R0_en = R0_en & R0_addr_sel == 8'h5f;
  assign mem_95_1_W0_addr = W0_addr[25:0];
  assign mem_95_1_W0_clk = W0_clk;
  assign mem_95_1_W0_data = W0_data[15:8];
  assign mem_95_1_W0_en = W0_en & W0_addr_sel == 8'h5f;
  assign mem_95_1_W0_mask = W0_mask[1];
  assign mem_95_2_R0_addr = R0_addr[25:0];
  assign mem_95_2_R0_clk = R0_clk;
  assign mem_95_2_R0_en = R0_en & R0_addr_sel == 8'h5f;
  assign mem_95_2_W0_addr = W0_addr[25:0];
  assign mem_95_2_W0_clk = W0_clk;
  assign mem_95_2_W0_data = W0_data[23:16];
  assign mem_95_2_W0_en = W0_en & W0_addr_sel == 8'h5f;
  assign mem_95_2_W0_mask = W0_mask[2];
  assign mem_95_3_R0_addr = R0_addr[25:0];
  assign mem_95_3_R0_clk = R0_clk;
  assign mem_95_3_R0_en = R0_en & R0_addr_sel == 8'h5f;
  assign mem_95_3_W0_addr = W0_addr[25:0];
  assign mem_95_3_W0_clk = W0_clk;
  assign mem_95_3_W0_data = W0_data[31:24];
  assign mem_95_3_W0_en = W0_en & W0_addr_sel == 8'h5f;
  assign mem_95_3_W0_mask = W0_mask[3];
  assign mem_95_4_R0_addr = R0_addr[25:0];
  assign mem_95_4_R0_clk = R0_clk;
  assign mem_95_4_R0_en = R0_en & R0_addr_sel == 8'h5f;
  assign mem_95_4_W0_addr = W0_addr[25:0];
  assign mem_95_4_W0_clk = W0_clk;
  assign mem_95_4_W0_data = W0_data[39:32];
  assign mem_95_4_W0_en = W0_en & W0_addr_sel == 8'h5f;
  assign mem_95_4_W0_mask = W0_mask[4];
  assign mem_95_5_R0_addr = R0_addr[25:0];
  assign mem_95_5_R0_clk = R0_clk;
  assign mem_95_5_R0_en = R0_en & R0_addr_sel == 8'h5f;
  assign mem_95_5_W0_addr = W0_addr[25:0];
  assign mem_95_5_W0_clk = W0_clk;
  assign mem_95_5_W0_data = W0_data[47:40];
  assign mem_95_5_W0_en = W0_en & W0_addr_sel == 8'h5f;
  assign mem_95_5_W0_mask = W0_mask[5];
  assign mem_95_6_R0_addr = R0_addr[25:0];
  assign mem_95_6_R0_clk = R0_clk;
  assign mem_95_6_R0_en = R0_en & R0_addr_sel == 8'h5f;
  assign mem_95_6_W0_addr = W0_addr[25:0];
  assign mem_95_6_W0_clk = W0_clk;
  assign mem_95_6_W0_data = W0_data[55:48];
  assign mem_95_6_W0_en = W0_en & W0_addr_sel == 8'h5f;
  assign mem_95_6_W0_mask = W0_mask[6];
  assign mem_95_7_R0_addr = R0_addr[25:0];
  assign mem_95_7_R0_clk = R0_clk;
  assign mem_95_7_R0_en = R0_en & R0_addr_sel == 8'h5f;
  assign mem_95_7_W0_addr = W0_addr[25:0];
  assign mem_95_7_W0_clk = W0_clk;
  assign mem_95_7_W0_data = W0_data[63:56];
  assign mem_95_7_W0_en = W0_en & W0_addr_sel == 8'h5f;
  assign mem_95_7_W0_mask = W0_mask[7];
  assign mem_96_0_R0_addr = R0_addr[25:0];
  assign mem_96_0_R0_clk = R0_clk;
  assign mem_96_0_R0_en = R0_en & R0_addr_sel == 8'h60;
  assign mem_96_0_W0_addr = W0_addr[25:0];
  assign mem_96_0_W0_clk = W0_clk;
  assign mem_96_0_W0_data = W0_data[7:0];
  assign mem_96_0_W0_en = W0_en & W0_addr_sel == 8'h60;
  assign mem_96_0_W0_mask = W0_mask[0];
  assign mem_96_1_R0_addr = R0_addr[25:0];
  assign mem_96_1_R0_clk = R0_clk;
  assign mem_96_1_R0_en = R0_en & R0_addr_sel == 8'h60;
  assign mem_96_1_W0_addr = W0_addr[25:0];
  assign mem_96_1_W0_clk = W0_clk;
  assign mem_96_1_W0_data = W0_data[15:8];
  assign mem_96_1_W0_en = W0_en & W0_addr_sel == 8'h60;
  assign mem_96_1_W0_mask = W0_mask[1];
  assign mem_96_2_R0_addr = R0_addr[25:0];
  assign mem_96_2_R0_clk = R0_clk;
  assign mem_96_2_R0_en = R0_en & R0_addr_sel == 8'h60;
  assign mem_96_2_W0_addr = W0_addr[25:0];
  assign mem_96_2_W0_clk = W0_clk;
  assign mem_96_2_W0_data = W0_data[23:16];
  assign mem_96_2_W0_en = W0_en & W0_addr_sel == 8'h60;
  assign mem_96_2_W0_mask = W0_mask[2];
  assign mem_96_3_R0_addr = R0_addr[25:0];
  assign mem_96_3_R0_clk = R0_clk;
  assign mem_96_3_R0_en = R0_en & R0_addr_sel == 8'h60;
  assign mem_96_3_W0_addr = W0_addr[25:0];
  assign mem_96_3_W0_clk = W0_clk;
  assign mem_96_3_W0_data = W0_data[31:24];
  assign mem_96_3_W0_en = W0_en & W0_addr_sel == 8'h60;
  assign mem_96_3_W0_mask = W0_mask[3];
  assign mem_96_4_R0_addr = R0_addr[25:0];
  assign mem_96_4_R0_clk = R0_clk;
  assign mem_96_4_R0_en = R0_en & R0_addr_sel == 8'h60;
  assign mem_96_4_W0_addr = W0_addr[25:0];
  assign mem_96_4_W0_clk = W0_clk;
  assign mem_96_4_W0_data = W0_data[39:32];
  assign mem_96_4_W0_en = W0_en & W0_addr_sel == 8'h60;
  assign mem_96_4_W0_mask = W0_mask[4];
  assign mem_96_5_R0_addr = R0_addr[25:0];
  assign mem_96_5_R0_clk = R0_clk;
  assign mem_96_5_R0_en = R0_en & R0_addr_sel == 8'h60;
  assign mem_96_5_W0_addr = W0_addr[25:0];
  assign mem_96_5_W0_clk = W0_clk;
  assign mem_96_5_W0_data = W0_data[47:40];
  assign mem_96_5_W0_en = W0_en & W0_addr_sel == 8'h60;
  assign mem_96_5_W0_mask = W0_mask[5];
  assign mem_96_6_R0_addr = R0_addr[25:0];
  assign mem_96_6_R0_clk = R0_clk;
  assign mem_96_6_R0_en = R0_en & R0_addr_sel == 8'h60;
  assign mem_96_6_W0_addr = W0_addr[25:0];
  assign mem_96_6_W0_clk = W0_clk;
  assign mem_96_6_W0_data = W0_data[55:48];
  assign mem_96_6_W0_en = W0_en & W0_addr_sel == 8'h60;
  assign mem_96_6_W0_mask = W0_mask[6];
  assign mem_96_7_R0_addr = R0_addr[25:0];
  assign mem_96_7_R0_clk = R0_clk;
  assign mem_96_7_R0_en = R0_en & R0_addr_sel == 8'h60;
  assign mem_96_7_W0_addr = W0_addr[25:0];
  assign mem_96_7_W0_clk = W0_clk;
  assign mem_96_7_W0_data = W0_data[63:56];
  assign mem_96_7_W0_en = W0_en & W0_addr_sel == 8'h60;
  assign mem_96_7_W0_mask = W0_mask[7];
  assign mem_97_0_R0_addr = R0_addr[25:0];
  assign mem_97_0_R0_clk = R0_clk;
  assign mem_97_0_R0_en = R0_en & R0_addr_sel == 8'h61;
  assign mem_97_0_W0_addr = W0_addr[25:0];
  assign mem_97_0_W0_clk = W0_clk;
  assign mem_97_0_W0_data = W0_data[7:0];
  assign mem_97_0_W0_en = W0_en & W0_addr_sel == 8'h61;
  assign mem_97_0_W0_mask = W0_mask[0];
  assign mem_97_1_R0_addr = R0_addr[25:0];
  assign mem_97_1_R0_clk = R0_clk;
  assign mem_97_1_R0_en = R0_en & R0_addr_sel == 8'h61;
  assign mem_97_1_W0_addr = W0_addr[25:0];
  assign mem_97_1_W0_clk = W0_clk;
  assign mem_97_1_W0_data = W0_data[15:8];
  assign mem_97_1_W0_en = W0_en & W0_addr_sel == 8'h61;
  assign mem_97_1_W0_mask = W0_mask[1];
  assign mem_97_2_R0_addr = R0_addr[25:0];
  assign mem_97_2_R0_clk = R0_clk;
  assign mem_97_2_R0_en = R0_en & R0_addr_sel == 8'h61;
  assign mem_97_2_W0_addr = W0_addr[25:0];
  assign mem_97_2_W0_clk = W0_clk;
  assign mem_97_2_W0_data = W0_data[23:16];
  assign mem_97_2_W0_en = W0_en & W0_addr_sel == 8'h61;
  assign mem_97_2_W0_mask = W0_mask[2];
  assign mem_97_3_R0_addr = R0_addr[25:0];
  assign mem_97_3_R0_clk = R0_clk;
  assign mem_97_3_R0_en = R0_en & R0_addr_sel == 8'h61;
  assign mem_97_3_W0_addr = W0_addr[25:0];
  assign mem_97_3_W0_clk = W0_clk;
  assign mem_97_3_W0_data = W0_data[31:24];
  assign mem_97_3_W0_en = W0_en & W0_addr_sel == 8'h61;
  assign mem_97_3_W0_mask = W0_mask[3];
  assign mem_97_4_R0_addr = R0_addr[25:0];
  assign mem_97_4_R0_clk = R0_clk;
  assign mem_97_4_R0_en = R0_en & R0_addr_sel == 8'h61;
  assign mem_97_4_W0_addr = W0_addr[25:0];
  assign mem_97_4_W0_clk = W0_clk;
  assign mem_97_4_W0_data = W0_data[39:32];
  assign mem_97_4_W0_en = W0_en & W0_addr_sel == 8'h61;
  assign mem_97_4_W0_mask = W0_mask[4];
  assign mem_97_5_R0_addr = R0_addr[25:0];
  assign mem_97_5_R0_clk = R0_clk;
  assign mem_97_5_R0_en = R0_en & R0_addr_sel == 8'h61;
  assign mem_97_5_W0_addr = W0_addr[25:0];
  assign mem_97_5_W0_clk = W0_clk;
  assign mem_97_5_W0_data = W0_data[47:40];
  assign mem_97_5_W0_en = W0_en & W0_addr_sel == 8'h61;
  assign mem_97_5_W0_mask = W0_mask[5];
  assign mem_97_6_R0_addr = R0_addr[25:0];
  assign mem_97_6_R0_clk = R0_clk;
  assign mem_97_6_R0_en = R0_en & R0_addr_sel == 8'h61;
  assign mem_97_6_W0_addr = W0_addr[25:0];
  assign mem_97_6_W0_clk = W0_clk;
  assign mem_97_6_W0_data = W0_data[55:48];
  assign mem_97_6_W0_en = W0_en & W0_addr_sel == 8'h61;
  assign mem_97_6_W0_mask = W0_mask[6];
  assign mem_97_7_R0_addr = R0_addr[25:0];
  assign mem_97_7_R0_clk = R0_clk;
  assign mem_97_7_R0_en = R0_en & R0_addr_sel == 8'h61;
  assign mem_97_7_W0_addr = W0_addr[25:0];
  assign mem_97_7_W0_clk = W0_clk;
  assign mem_97_7_W0_data = W0_data[63:56];
  assign mem_97_7_W0_en = W0_en & W0_addr_sel == 8'h61;
  assign mem_97_7_W0_mask = W0_mask[7];
  assign mem_98_0_R0_addr = R0_addr[25:0];
  assign mem_98_0_R0_clk = R0_clk;
  assign mem_98_0_R0_en = R0_en & R0_addr_sel == 8'h62;
  assign mem_98_0_W0_addr = W0_addr[25:0];
  assign mem_98_0_W0_clk = W0_clk;
  assign mem_98_0_W0_data = W0_data[7:0];
  assign mem_98_0_W0_en = W0_en & W0_addr_sel == 8'h62;
  assign mem_98_0_W0_mask = W0_mask[0];
  assign mem_98_1_R0_addr = R0_addr[25:0];
  assign mem_98_1_R0_clk = R0_clk;
  assign mem_98_1_R0_en = R0_en & R0_addr_sel == 8'h62;
  assign mem_98_1_W0_addr = W0_addr[25:0];
  assign mem_98_1_W0_clk = W0_clk;
  assign mem_98_1_W0_data = W0_data[15:8];
  assign mem_98_1_W0_en = W0_en & W0_addr_sel == 8'h62;
  assign mem_98_1_W0_mask = W0_mask[1];
  assign mem_98_2_R0_addr = R0_addr[25:0];
  assign mem_98_2_R0_clk = R0_clk;
  assign mem_98_2_R0_en = R0_en & R0_addr_sel == 8'h62;
  assign mem_98_2_W0_addr = W0_addr[25:0];
  assign mem_98_2_W0_clk = W0_clk;
  assign mem_98_2_W0_data = W0_data[23:16];
  assign mem_98_2_W0_en = W0_en & W0_addr_sel == 8'h62;
  assign mem_98_2_W0_mask = W0_mask[2];
  assign mem_98_3_R0_addr = R0_addr[25:0];
  assign mem_98_3_R0_clk = R0_clk;
  assign mem_98_3_R0_en = R0_en & R0_addr_sel == 8'h62;
  assign mem_98_3_W0_addr = W0_addr[25:0];
  assign mem_98_3_W0_clk = W0_clk;
  assign mem_98_3_W0_data = W0_data[31:24];
  assign mem_98_3_W0_en = W0_en & W0_addr_sel == 8'h62;
  assign mem_98_3_W0_mask = W0_mask[3];
  assign mem_98_4_R0_addr = R0_addr[25:0];
  assign mem_98_4_R0_clk = R0_clk;
  assign mem_98_4_R0_en = R0_en & R0_addr_sel == 8'h62;
  assign mem_98_4_W0_addr = W0_addr[25:0];
  assign mem_98_4_W0_clk = W0_clk;
  assign mem_98_4_W0_data = W0_data[39:32];
  assign mem_98_4_W0_en = W0_en & W0_addr_sel == 8'h62;
  assign mem_98_4_W0_mask = W0_mask[4];
  assign mem_98_5_R0_addr = R0_addr[25:0];
  assign mem_98_5_R0_clk = R0_clk;
  assign mem_98_5_R0_en = R0_en & R0_addr_sel == 8'h62;
  assign mem_98_5_W0_addr = W0_addr[25:0];
  assign mem_98_5_W0_clk = W0_clk;
  assign mem_98_5_W0_data = W0_data[47:40];
  assign mem_98_5_W0_en = W0_en & W0_addr_sel == 8'h62;
  assign mem_98_5_W0_mask = W0_mask[5];
  assign mem_98_6_R0_addr = R0_addr[25:0];
  assign mem_98_6_R0_clk = R0_clk;
  assign mem_98_6_R0_en = R0_en & R0_addr_sel == 8'h62;
  assign mem_98_6_W0_addr = W0_addr[25:0];
  assign mem_98_6_W0_clk = W0_clk;
  assign mem_98_6_W0_data = W0_data[55:48];
  assign mem_98_6_W0_en = W0_en & W0_addr_sel == 8'h62;
  assign mem_98_6_W0_mask = W0_mask[6];
  assign mem_98_7_R0_addr = R0_addr[25:0];
  assign mem_98_7_R0_clk = R0_clk;
  assign mem_98_7_R0_en = R0_en & R0_addr_sel == 8'h62;
  assign mem_98_7_W0_addr = W0_addr[25:0];
  assign mem_98_7_W0_clk = W0_clk;
  assign mem_98_7_W0_data = W0_data[63:56];
  assign mem_98_7_W0_en = W0_en & W0_addr_sel == 8'h62;
  assign mem_98_7_W0_mask = W0_mask[7];
  assign mem_99_0_R0_addr = R0_addr[25:0];
  assign mem_99_0_R0_clk = R0_clk;
  assign mem_99_0_R0_en = R0_en & R0_addr_sel == 8'h63;
  assign mem_99_0_W0_addr = W0_addr[25:0];
  assign mem_99_0_W0_clk = W0_clk;
  assign mem_99_0_W0_data = W0_data[7:0];
  assign mem_99_0_W0_en = W0_en & W0_addr_sel == 8'h63;
  assign mem_99_0_W0_mask = W0_mask[0];
  assign mem_99_1_R0_addr = R0_addr[25:0];
  assign mem_99_1_R0_clk = R0_clk;
  assign mem_99_1_R0_en = R0_en & R0_addr_sel == 8'h63;
  assign mem_99_1_W0_addr = W0_addr[25:0];
  assign mem_99_1_W0_clk = W0_clk;
  assign mem_99_1_W0_data = W0_data[15:8];
  assign mem_99_1_W0_en = W0_en & W0_addr_sel == 8'h63;
  assign mem_99_1_W0_mask = W0_mask[1];
  assign mem_99_2_R0_addr = R0_addr[25:0];
  assign mem_99_2_R0_clk = R0_clk;
  assign mem_99_2_R0_en = R0_en & R0_addr_sel == 8'h63;
  assign mem_99_2_W0_addr = W0_addr[25:0];
  assign mem_99_2_W0_clk = W0_clk;
  assign mem_99_2_W0_data = W0_data[23:16];
  assign mem_99_2_W0_en = W0_en & W0_addr_sel == 8'h63;
  assign mem_99_2_W0_mask = W0_mask[2];
  assign mem_99_3_R0_addr = R0_addr[25:0];
  assign mem_99_3_R0_clk = R0_clk;
  assign mem_99_3_R0_en = R0_en & R0_addr_sel == 8'h63;
  assign mem_99_3_W0_addr = W0_addr[25:0];
  assign mem_99_3_W0_clk = W0_clk;
  assign mem_99_3_W0_data = W0_data[31:24];
  assign mem_99_3_W0_en = W0_en & W0_addr_sel == 8'h63;
  assign mem_99_3_W0_mask = W0_mask[3];
  assign mem_99_4_R0_addr = R0_addr[25:0];
  assign mem_99_4_R0_clk = R0_clk;
  assign mem_99_4_R0_en = R0_en & R0_addr_sel == 8'h63;
  assign mem_99_4_W0_addr = W0_addr[25:0];
  assign mem_99_4_W0_clk = W0_clk;
  assign mem_99_4_W0_data = W0_data[39:32];
  assign mem_99_4_W0_en = W0_en & W0_addr_sel == 8'h63;
  assign mem_99_4_W0_mask = W0_mask[4];
  assign mem_99_5_R0_addr = R0_addr[25:0];
  assign mem_99_5_R0_clk = R0_clk;
  assign mem_99_5_R0_en = R0_en & R0_addr_sel == 8'h63;
  assign mem_99_5_W0_addr = W0_addr[25:0];
  assign mem_99_5_W0_clk = W0_clk;
  assign mem_99_5_W0_data = W0_data[47:40];
  assign mem_99_5_W0_en = W0_en & W0_addr_sel == 8'h63;
  assign mem_99_5_W0_mask = W0_mask[5];
  assign mem_99_6_R0_addr = R0_addr[25:0];
  assign mem_99_6_R0_clk = R0_clk;
  assign mem_99_6_R0_en = R0_en & R0_addr_sel == 8'h63;
  assign mem_99_6_W0_addr = W0_addr[25:0];
  assign mem_99_6_W0_clk = W0_clk;
  assign mem_99_6_W0_data = W0_data[55:48];
  assign mem_99_6_W0_en = W0_en & W0_addr_sel == 8'h63;
  assign mem_99_6_W0_mask = W0_mask[6];
  assign mem_99_7_R0_addr = R0_addr[25:0];
  assign mem_99_7_R0_clk = R0_clk;
  assign mem_99_7_R0_en = R0_en & R0_addr_sel == 8'h63;
  assign mem_99_7_W0_addr = W0_addr[25:0];
  assign mem_99_7_W0_clk = W0_clk;
  assign mem_99_7_W0_data = W0_data[63:56];
  assign mem_99_7_W0_en = W0_en & W0_addr_sel == 8'h63;
  assign mem_99_7_W0_mask = W0_mask[7];
  assign mem_100_0_R0_addr = R0_addr[25:0];
  assign mem_100_0_R0_clk = R0_clk;
  assign mem_100_0_R0_en = R0_en & R0_addr_sel == 8'h64;
  assign mem_100_0_W0_addr = W0_addr[25:0];
  assign mem_100_0_W0_clk = W0_clk;
  assign mem_100_0_W0_data = W0_data[7:0];
  assign mem_100_0_W0_en = W0_en & W0_addr_sel == 8'h64;
  assign mem_100_0_W0_mask = W0_mask[0];
  assign mem_100_1_R0_addr = R0_addr[25:0];
  assign mem_100_1_R0_clk = R0_clk;
  assign mem_100_1_R0_en = R0_en & R0_addr_sel == 8'h64;
  assign mem_100_1_W0_addr = W0_addr[25:0];
  assign mem_100_1_W0_clk = W0_clk;
  assign mem_100_1_W0_data = W0_data[15:8];
  assign mem_100_1_W0_en = W0_en & W0_addr_sel == 8'h64;
  assign mem_100_1_W0_mask = W0_mask[1];
  assign mem_100_2_R0_addr = R0_addr[25:0];
  assign mem_100_2_R0_clk = R0_clk;
  assign mem_100_2_R0_en = R0_en & R0_addr_sel == 8'h64;
  assign mem_100_2_W0_addr = W0_addr[25:0];
  assign mem_100_2_W0_clk = W0_clk;
  assign mem_100_2_W0_data = W0_data[23:16];
  assign mem_100_2_W0_en = W0_en & W0_addr_sel == 8'h64;
  assign mem_100_2_W0_mask = W0_mask[2];
  assign mem_100_3_R0_addr = R0_addr[25:0];
  assign mem_100_3_R0_clk = R0_clk;
  assign mem_100_3_R0_en = R0_en & R0_addr_sel == 8'h64;
  assign mem_100_3_W0_addr = W0_addr[25:0];
  assign mem_100_3_W0_clk = W0_clk;
  assign mem_100_3_W0_data = W0_data[31:24];
  assign mem_100_3_W0_en = W0_en & W0_addr_sel == 8'h64;
  assign mem_100_3_W0_mask = W0_mask[3];
  assign mem_100_4_R0_addr = R0_addr[25:0];
  assign mem_100_4_R0_clk = R0_clk;
  assign mem_100_4_R0_en = R0_en & R0_addr_sel == 8'h64;
  assign mem_100_4_W0_addr = W0_addr[25:0];
  assign mem_100_4_W0_clk = W0_clk;
  assign mem_100_4_W0_data = W0_data[39:32];
  assign mem_100_4_W0_en = W0_en & W0_addr_sel == 8'h64;
  assign mem_100_4_W0_mask = W0_mask[4];
  assign mem_100_5_R0_addr = R0_addr[25:0];
  assign mem_100_5_R0_clk = R0_clk;
  assign mem_100_5_R0_en = R0_en & R0_addr_sel == 8'h64;
  assign mem_100_5_W0_addr = W0_addr[25:0];
  assign mem_100_5_W0_clk = W0_clk;
  assign mem_100_5_W0_data = W0_data[47:40];
  assign mem_100_5_W0_en = W0_en & W0_addr_sel == 8'h64;
  assign mem_100_5_W0_mask = W0_mask[5];
  assign mem_100_6_R0_addr = R0_addr[25:0];
  assign mem_100_6_R0_clk = R0_clk;
  assign mem_100_6_R0_en = R0_en & R0_addr_sel == 8'h64;
  assign mem_100_6_W0_addr = W0_addr[25:0];
  assign mem_100_6_W0_clk = W0_clk;
  assign mem_100_6_W0_data = W0_data[55:48];
  assign mem_100_6_W0_en = W0_en & W0_addr_sel == 8'h64;
  assign mem_100_6_W0_mask = W0_mask[6];
  assign mem_100_7_R0_addr = R0_addr[25:0];
  assign mem_100_7_R0_clk = R0_clk;
  assign mem_100_7_R0_en = R0_en & R0_addr_sel == 8'h64;
  assign mem_100_7_W0_addr = W0_addr[25:0];
  assign mem_100_7_W0_clk = W0_clk;
  assign mem_100_7_W0_data = W0_data[63:56];
  assign mem_100_7_W0_en = W0_en & W0_addr_sel == 8'h64;
  assign mem_100_7_W0_mask = W0_mask[7];
  assign mem_101_0_R0_addr = R0_addr[25:0];
  assign mem_101_0_R0_clk = R0_clk;
  assign mem_101_0_R0_en = R0_en & R0_addr_sel == 8'h65;
  assign mem_101_0_W0_addr = W0_addr[25:0];
  assign mem_101_0_W0_clk = W0_clk;
  assign mem_101_0_W0_data = W0_data[7:0];
  assign mem_101_0_W0_en = W0_en & W0_addr_sel == 8'h65;
  assign mem_101_0_W0_mask = W0_mask[0];
  assign mem_101_1_R0_addr = R0_addr[25:0];
  assign mem_101_1_R0_clk = R0_clk;
  assign mem_101_1_R0_en = R0_en & R0_addr_sel == 8'h65;
  assign mem_101_1_W0_addr = W0_addr[25:0];
  assign mem_101_1_W0_clk = W0_clk;
  assign mem_101_1_W0_data = W0_data[15:8];
  assign mem_101_1_W0_en = W0_en & W0_addr_sel == 8'h65;
  assign mem_101_1_W0_mask = W0_mask[1];
  assign mem_101_2_R0_addr = R0_addr[25:0];
  assign mem_101_2_R0_clk = R0_clk;
  assign mem_101_2_R0_en = R0_en & R0_addr_sel == 8'h65;
  assign mem_101_2_W0_addr = W0_addr[25:0];
  assign mem_101_2_W0_clk = W0_clk;
  assign mem_101_2_W0_data = W0_data[23:16];
  assign mem_101_2_W0_en = W0_en & W0_addr_sel == 8'h65;
  assign mem_101_2_W0_mask = W0_mask[2];
  assign mem_101_3_R0_addr = R0_addr[25:0];
  assign mem_101_3_R0_clk = R0_clk;
  assign mem_101_3_R0_en = R0_en & R0_addr_sel == 8'h65;
  assign mem_101_3_W0_addr = W0_addr[25:0];
  assign mem_101_3_W0_clk = W0_clk;
  assign mem_101_3_W0_data = W0_data[31:24];
  assign mem_101_3_W0_en = W0_en & W0_addr_sel == 8'h65;
  assign mem_101_3_W0_mask = W0_mask[3];
  assign mem_101_4_R0_addr = R0_addr[25:0];
  assign mem_101_4_R0_clk = R0_clk;
  assign mem_101_4_R0_en = R0_en & R0_addr_sel == 8'h65;
  assign mem_101_4_W0_addr = W0_addr[25:0];
  assign mem_101_4_W0_clk = W0_clk;
  assign mem_101_4_W0_data = W0_data[39:32];
  assign mem_101_4_W0_en = W0_en & W0_addr_sel == 8'h65;
  assign mem_101_4_W0_mask = W0_mask[4];
  assign mem_101_5_R0_addr = R0_addr[25:0];
  assign mem_101_5_R0_clk = R0_clk;
  assign mem_101_5_R0_en = R0_en & R0_addr_sel == 8'h65;
  assign mem_101_5_W0_addr = W0_addr[25:0];
  assign mem_101_5_W0_clk = W0_clk;
  assign mem_101_5_W0_data = W0_data[47:40];
  assign mem_101_5_W0_en = W0_en & W0_addr_sel == 8'h65;
  assign mem_101_5_W0_mask = W0_mask[5];
  assign mem_101_6_R0_addr = R0_addr[25:0];
  assign mem_101_6_R0_clk = R0_clk;
  assign mem_101_6_R0_en = R0_en & R0_addr_sel == 8'h65;
  assign mem_101_6_W0_addr = W0_addr[25:0];
  assign mem_101_6_W0_clk = W0_clk;
  assign mem_101_6_W0_data = W0_data[55:48];
  assign mem_101_6_W0_en = W0_en & W0_addr_sel == 8'h65;
  assign mem_101_6_W0_mask = W0_mask[6];
  assign mem_101_7_R0_addr = R0_addr[25:0];
  assign mem_101_7_R0_clk = R0_clk;
  assign mem_101_7_R0_en = R0_en & R0_addr_sel == 8'h65;
  assign mem_101_7_W0_addr = W0_addr[25:0];
  assign mem_101_7_W0_clk = W0_clk;
  assign mem_101_7_W0_data = W0_data[63:56];
  assign mem_101_7_W0_en = W0_en & W0_addr_sel == 8'h65;
  assign mem_101_7_W0_mask = W0_mask[7];
  assign mem_102_0_R0_addr = R0_addr[25:0];
  assign mem_102_0_R0_clk = R0_clk;
  assign mem_102_0_R0_en = R0_en & R0_addr_sel == 8'h66;
  assign mem_102_0_W0_addr = W0_addr[25:0];
  assign mem_102_0_W0_clk = W0_clk;
  assign mem_102_0_W0_data = W0_data[7:0];
  assign mem_102_0_W0_en = W0_en & W0_addr_sel == 8'h66;
  assign mem_102_0_W0_mask = W0_mask[0];
  assign mem_102_1_R0_addr = R0_addr[25:0];
  assign mem_102_1_R0_clk = R0_clk;
  assign mem_102_1_R0_en = R0_en & R0_addr_sel == 8'h66;
  assign mem_102_1_W0_addr = W0_addr[25:0];
  assign mem_102_1_W0_clk = W0_clk;
  assign mem_102_1_W0_data = W0_data[15:8];
  assign mem_102_1_W0_en = W0_en & W0_addr_sel == 8'h66;
  assign mem_102_1_W0_mask = W0_mask[1];
  assign mem_102_2_R0_addr = R0_addr[25:0];
  assign mem_102_2_R0_clk = R0_clk;
  assign mem_102_2_R0_en = R0_en & R0_addr_sel == 8'h66;
  assign mem_102_2_W0_addr = W0_addr[25:0];
  assign mem_102_2_W0_clk = W0_clk;
  assign mem_102_2_W0_data = W0_data[23:16];
  assign mem_102_2_W0_en = W0_en & W0_addr_sel == 8'h66;
  assign mem_102_2_W0_mask = W0_mask[2];
  assign mem_102_3_R0_addr = R0_addr[25:0];
  assign mem_102_3_R0_clk = R0_clk;
  assign mem_102_3_R0_en = R0_en & R0_addr_sel == 8'h66;
  assign mem_102_3_W0_addr = W0_addr[25:0];
  assign mem_102_3_W0_clk = W0_clk;
  assign mem_102_3_W0_data = W0_data[31:24];
  assign mem_102_3_W0_en = W0_en & W0_addr_sel == 8'h66;
  assign mem_102_3_W0_mask = W0_mask[3];
  assign mem_102_4_R0_addr = R0_addr[25:0];
  assign mem_102_4_R0_clk = R0_clk;
  assign mem_102_4_R0_en = R0_en & R0_addr_sel == 8'h66;
  assign mem_102_4_W0_addr = W0_addr[25:0];
  assign mem_102_4_W0_clk = W0_clk;
  assign mem_102_4_W0_data = W0_data[39:32];
  assign mem_102_4_W0_en = W0_en & W0_addr_sel == 8'h66;
  assign mem_102_4_W0_mask = W0_mask[4];
  assign mem_102_5_R0_addr = R0_addr[25:0];
  assign mem_102_5_R0_clk = R0_clk;
  assign mem_102_5_R0_en = R0_en & R0_addr_sel == 8'h66;
  assign mem_102_5_W0_addr = W0_addr[25:0];
  assign mem_102_5_W0_clk = W0_clk;
  assign mem_102_5_W0_data = W0_data[47:40];
  assign mem_102_5_W0_en = W0_en & W0_addr_sel == 8'h66;
  assign mem_102_5_W0_mask = W0_mask[5];
  assign mem_102_6_R0_addr = R0_addr[25:0];
  assign mem_102_6_R0_clk = R0_clk;
  assign mem_102_6_R0_en = R0_en & R0_addr_sel == 8'h66;
  assign mem_102_6_W0_addr = W0_addr[25:0];
  assign mem_102_6_W0_clk = W0_clk;
  assign mem_102_6_W0_data = W0_data[55:48];
  assign mem_102_6_W0_en = W0_en & W0_addr_sel == 8'h66;
  assign mem_102_6_W0_mask = W0_mask[6];
  assign mem_102_7_R0_addr = R0_addr[25:0];
  assign mem_102_7_R0_clk = R0_clk;
  assign mem_102_7_R0_en = R0_en & R0_addr_sel == 8'h66;
  assign mem_102_7_W0_addr = W0_addr[25:0];
  assign mem_102_7_W0_clk = W0_clk;
  assign mem_102_7_W0_data = W0_data[63:56];
  assign mem_102_7_W0_en = W0_en & W0_addr_sel == 8'h66;
  assign mem_102_7_W0_mask = W0_mask[7];
  assign mem_103_0_R0_addr = R0_addr[25:0];
  assign mem_103_0_R0_clk = R0_clk;
  assign mem_103_0_R0_en = R0_en & R0_addr_sel == 8'h67;
  assign mem_103_0_W0_addr = W0_addr[25:0];
  assign mem_103_0_W0_clk = W0_clk;
  assign mem_103_0_W0_data = W0_data[7:0];
  assign mem_103_0_W0_en = W0_en & W0_addr_sel == 8'h67;
  assign mem_103_0_W0_mask = W0_mask[0];
  assign mem_103_1_R0_addr = R0_addr[25:0];
  assign mem_103_1_R0_clk = R0_clk;
  assign mem_103_1_R0_en = R0_en & R0_addr_sel == 8'h67;
  assign mem_103_1_W0_addr = W0_addr[25:0];
  assign mem_103_1_W0_clk = W0_clk;
  assign mem_103_1_W0_data = W0_data[15:8];
  assign mem_103_1_W0_en = W0_en & W0_addr_sel == 8'h67;
  assign mem_103_1_W0_mask = W0_mask[1];
  assign mem_103_2_R0_addr = R0_addr[25:0];
  assign mem_103_2_R0_clk = R0_clk;
  assign mem_103_2_R0_en = R0_en & R0_addr_sel == 8'h67;
  assign mem_103_2_W0_addr = W0_addr[25:0];
  assign mem_103_2_W0_clk = W0_clk;
  assign mem_103_2_W0_data = W0_data[23:16];
  assign mem_103_2_W0_en = W0_en & W0_addr_sel == 8'h67;
  assign mem_103_2_W0_mask = W0_mask[2];
  assign mem_103_3_R0_addr = R0_addr[25:0];
  assign mem_103_3_R0_clk = R0_clk;
  assign mem_103_3_R0_en = R0_en & R0_addr_sel == 8'h67;
  assign mem_103_3_W0_addr = W0_addr[25:0];
  assign mem_103_3_W0_clk = W0_clk;
  assign mem_103_3_W0_data = W0_data[31:24];
  assign mem_103_3_W0_en = W0_en & W0_addr_sel == 8'h67;
  assign mem_103_3_W0_mask = W0_mask[3];
  assign mem_103_4_R0_addr = R0_addr[25:0];
  assign mem_103_4_R0_clk = R0_clk;
  assign mem_103_4_R0_en = R0_en & R0_addr_sel == 8'h67;
  assign mem_103_4_W0_addr = W0_addr[25:0];
  assign mem_103_4_W0_clk = W0_clk;
  assign mem_103_4_W0_data = W0_data[39:32];
  assign mem_103_4_W0_en = W0_en & W0_addr_sel == 8'h67;
  assign mem_103_4_W0_mask = W0_mask[4];
  assign mem_103_5_R0_addr = R0_addr[25:0];
  assign mem_103_5_R0_clk = R0_clk;
  assign mem_103_5_R0_en = R0_en & R0_addr_sel == 8'h67;
  assign mem_103_5_W0_addr = W0_addr[25:0];
  assign mem_103_5_W0_clk = W0_clk;
  assign mem_103_5_W0_data = W0_data[47:40];
  assign mem_103_5_W0_en = W0_en & W0_addr_sel == 8'h67;
  assign mem_103_5_W0_mask = W0_mask[5];
  assign mem_103_6_R0_addr = R0_addr[25:0];
  assign mem_103_6_R0_clk = R0_clk;
  assign mem_103_6_R0_en = R0_en & R0_addr_sel == 8'h67;
  assign mem_103_6_W0_addr = W0_addr[25:0];
  assign mem_103_6_W0_clk = W0_clk;
  assign mem_103_6_W0_data = W0_data[55:48];
  assign mem_103_6_W0_en = W0_en & W0_addr_sel == 8'h67;
  assign mem_103_6_W0_mask = W0_mask[6];
  assign mem_103_7_R0_addr = R0_addr[25:0];
  assign mem_103_7_R0_clk = R0_clk;
  assign mem_103_7_R0_en = R0_en & R0_addr_sel == 8'h67;
  assign mem_103_7_W0_addr = W0_addr[25:0];
  assign mem_103_7_W0_clk = W0_clk;
  assign mem_103_7_W0_data = W0_data[63:56];
  assign mem_103_7_W0_en = W0_en & W0_addr_sel == 8'h67;
  assign mem_103_7_W0_mask = W0_mask[7];
  assign mem_104_0_R0_addr = R0_addr[25:0];
  assign mem_104_0_R0_clk = R0_clk;
  assign mem_104_0_R0_en = R0_en & R0_addr_sel == 8'h68;
  assign mem_104_0_W0_addr = W0_addr[25:0];
  assign mem_104_0_W0_clk = W0_clk;
  assign mem_104_0_W0_data = W0_data[7:0];
  assign mem_104_0_W0_en = W0_en & W0_addr_sel == 8'h68;
  assign mem_104_0_W0_mask = W0_mask[0];
  assign mem_104_1_R0_addr = R0_addr[25:0];
  assign mem_104_1_R0_clk = R0_clk;
  assign mem_104_1_R0_en = R0_en & R0_addr_sel == 8'h68;
  assign mem_104_1_W0_addr = W0_addr[25:0];
  assign mem_104_1_W0_clk = W0_clk;
  assign mem_104_1_W0_data = W0_data[15:8];
  assign mem_104_1_W0_en = W0_en & W0_addr_sel == 8'h68;
  assign mem_104_1_W0_mask = W0_mask[1];
  assign mem_104_2_R0_addr = R0_addr[25:0];
  assign mem_104_2_R0_clk = R0_clk;
  assign mem_104_2_R0_en = R0_en & R0_addr_sel == 8'h68;
  assign mem_104_2_W0_addr = W0_addr[25:0];
  assign mem_104_2_W0_clk = W0_clk;
  assign mem_104_2_W0_data = W0_data[23:16];
  assign mem_104_2_W0_en = W0_en & W0_addr_sel == 8'h68;
  assign mem_104_2_W0_mask = W0_mask[2];
  assign mem_104_3_R0_addr = R0_addr[25:0];
  assign mem_104_3_R0_clk = R0_clk;
  assign mem_104_3_R0_en = R0_en & R0_addr_sel == 8'h68;
  assign mem_104_3_W0_addr = W0_addr[25:0];
  assign mem_104_3_W0_clk = W0_clk;
  assign mem_104_3_W0_data = W0_data[31:24];
  assign mem_104_3_W0_en = W0_en & W0_addr_sel == 8'h68;
  assign mem_104_3_W0_mask = W0_mask[3];
  assign mem_104_4_R0_addr = R0_addr[25:0];
  assign mem_104_4_R0_clk = R0_clk;
  assign mem_104_4_R0_en = R0_en & R0_addr_sel == 8'h68;
  assign mem_104_4_W0_addr = W0_addr[25:0];
  assign mem_104_4_W0_clk = W0_clk;
  assign mem_104_4_W0_data = W0_data[39:32];
  assign mem_104_4_W0_en = W0_en & W0_addr_sel == 8'h68;
  assign mem_104_4_W0_mask = W0_mask[4];
  assign mem_104_5_R0_addr = R0_addr[25:0];
  assign mem_104_5_R0_clk = R0_clk;
  assign mem_104_5_R0_en = R0_en & R0_addr_sel == 8'h68;
  assign mem_104_5_W0_addr = W0_addr[25:0];
  assign mem_104_5_W0_clk = W0_clk;
  assign mem_104_5_W0_data = W0_data[47:40];
  assign mem_104_5_W0_en = W0_en & W0_addr_sel == 8'h68;
  assign mem_104_5_W0_mask = W0_mask[5];
  assign mem_104_6_R0_addr = R0_addr[25:0];
  assign mem_104_6_R0_clk = R0_clk;
  assign mem_104_6_R0_en = R0_en & R0_addr_sel == 8'h68;
  assign mem_104_6_W0_addr = W0_addr[25:0];
  assign mem_104_6_W0_clk = W0_clk;
  assign mem_104_6_W0_data = W0_data[55:48];
  assign mem_104_6_W0_en = W0_en & W0_addr_sel == 8'h68;
  assign mem_104_6_W0_mask = W0_mask[6];
  assign mem_104_7_R0_addr = R0_addr[25:0];
  assign mem_104_7_R0_clk = R0_clk;
  assign mem_104_7_R0_en = R0_en & R0_addr_sel == 8'h68;
  assign mem_104_7_W0_addr = W0_addr[25:0];
  assign mem_104_7_W0_clk = W0_clk;
  assign mem_104_7_W0_data = W0_data[63:56];
  assign mem_104_7_W0_en = W0_en & W0_addr_sel == 8'h68;
  assign mem_104_7_W0_mask = W0_mask[7];
  assign mem_105_0_R0_addr = R0_addr[25:0];
  assign mem_105_0_R0_clk = R0_clk;
  assign mem_105_0_R0_en = R0_en & R0_addr_sel == 8'h69;
  assign mem_105_0_W0_addr = W0_addr[25:0];
  assign mem_105_0_W0_clk = W0_clk;
  assign mem_105_0_W0_data = W0_data[7:0];
  assign mem_105_0_W0_en = W0_en & W0_addr_sel == 8'h69;
  assign mem_105_0_W0_mask = W0_mask[0];
  assign mem_105_1_R0_addr = R0_addr[25:0];
  assign mem_105_1_R0_clk = R0_clk;
  assign mem_105_1_R0_en = R0_en & R0_addr_sel == 8'h69;
  assign mem_105_1_W0_addr = W0_addr[25:0];
  assign mem_105_1_W0_clk = W0_clk;
  assign mem_105_1_W0_data = W0_data[15:8];
  assign mem_105_1_W0_en = W0_en & W0_addr_sel == 8'h69;
  assign mem_105_1_W0_mask = W0_mask[1];
  assign mem_105_2_R0_addr = R0_addr[25:0];
  assign mem_105_2_R0_clk = R0_clk;
  assign mem_105_2_R0_en = R0_en & R0_addr_sel == 8'h69;
  assign mem_105_2_W0_addr = W0_addr[25:0];
  assign mem_105_2_W0_clk = W0_clk;
  assign mem_105_2_W0_data = W0_data[23:16];
  assign mem_105_2_W0_en = W0_en & W0_addr_sel == 8'h69;
  assign mem_105_2_W0_mask = W0_mask[2];
  assign mem_105_3_R0_addr = R0_addr[25:0];
  assign mem_105_3_R0_clk = R0_clk;
  assign mem_105_3_R0_en = R0_en & R0_addr_sel == 8'h69;
  assign mem_105_3_W0_addr = W0_addr[25:0];
  assign mem_105_3_W0_clk = W0_clk;
  assign mem_105_3_W0_data = W0_data[31:24];
  assign mem_105_3_W0_en = W0_en & W0_addr_sel == 8'h69;
  assign mem_105_3_W0_mask = W0_mask[3];
  assign mem_105_4_R0_addr = R0_addr[25:0];
  assign mem_105_4_R0_clk = R0_clk;
  assign mem_105_4_R0_en = R0_en & R0_addr_sel == 8'h69;
  assign mem_105_4_W0_addr = W0_addr[25:0];
  assign mem_105_4_W0_clk = W0_clk;
  assign mem_105_4_W0_data = W0_data[39:32];
  assign mem_105_4_W0_en = W0_en & W0_addr_sel == 8'h69;
  assign mem_105_4_W0_mask = W0_mask[4];
  assign mem_105_5_R0_addr = R0_addr[25:0];
  assign mem_105_5_R0_clk = R0_clk;
  assign mem_105_5_R0_en = R0_en & R0_addr_sel == 8'h69;
  assign mem_105_5_W0_addr = W0_addr[25:0];
  assign mem_105_5_W0_clk = W0_clk;
  assign mem_105_5_W0_data = W0_data[47:40];
  assign mem_105_5_W0_en = W0_en & W0_addr_sel == 8'h69;
  assign mem_105_5_W0_mask = W0_mask[5];
  assign mem_105_6_R0_addr = R0_addr[25:0];
  assign mem_105_6_R0_clk = R0_clk;
  assign mem_105_6_R0_en = R0_en & R0_addr_sel == 8'h69;
  assign mem_105_6_W0_addr = W0_addr[25:0];
  assign mem_105_6_W0_clk = W0_clk;
  assign mem_105_6_W0_data = W0_data[55:48];
  assign mem_105_6_W0_en = W0_en & W0_addr_sel == 8'h69;
  assign mem_105_6_W0_mask = W0_mask[6];
  assign mem_105_7_R0_addr = R0_addr[25:0];
  assign mem_105_7_R0_clk = R0_clk;
  assign mem_105_7_R0_en = R0_en & R0_addr_sel == 8'h69;
  assign mem_105_7_W0_addr = W0_addr[25:0];
  assign mem_105_7_W0_clk = W0_clk;
  assign mem_105_7_W0_data = W0_data[63:56];
  assign mem_105_7_W0_en = W0_en & W0_addr_sel == 8'h69;
  assign mem_105_7_W0_mask = W0_mask[7];
  assign mem_106_0_R0_addr = R0_addr[25:0];
  assign mem_106_0_R0_clk = R0_clk;
  assign mem_106_0_R0_en = R0_en & R0_addr_sel == 8'h6a;
  assign mem_106_0_W0_addr = W0_addr[25:0];
  assign mem_106_0_W0_clk = W0_clk;
  assign mem_106_0_W0_data = W0_data[7:0];
  assign mem_106_0_W0_en = W0_en & W0_addr_sel == 8'h6a;
  assign mem_106_0_W0_mask = W0_mask[0];
  assign mem_106_1_R0_addr = R0_addr[25:0];
  assign mem_106_1_R0_clk = R0_clk;
  assign mem_106_1_R0_en = R0_en & R0_addr_sel == 8'h6a;
  assign mem_106_1_W0_addr = W0_addr[25:0];
  assign mem_106_1_W0_clk = W0_clk;
  assign mem_106_1_W0_data = W0_data[15:8];
  assign mem_106_1_W0_en = W0_en & W0_addr_sel == 8'h6a;
  assign mem_106_1_W0_mask = W0_mask[1];
  assign mem_106_2_R0_addr = R0_addr[25:0];
  assign mem_106_2_R0_clk = R0_clk;
  assign mem_106_2_R0_en = R0_en & R0_addr_sel == 8'h6a;
  assign mem_106_2_W0_addr = W0_addr[25:0];
  assign mem_106_2_W0_clk = W0_clk;
  assign mem_106_2_W0_data = W0_data[23:16];
  assign mem_106_2_W0_en = W0_en & W0_addr_sel == 8'h6a;
  assign mem_106_2_W0_mask = W0_mask[2];
  assign mem_106_3_R0_addr = R0_addr[25:0];
  assign mem_106_3_R0_clk = R0_clk;
  assign mem_106_3_R0_en = R0_en & R0_addr_sel == 8'h6a;
  assign mem_106_3_W0_addr = W0_addr[25:0];
  assign mem_106_3_W0_clk = W0_clk;
  assign mem_106_3_W0_data = W0_data[31:24];
  assign mem_106_3_W0_en = W0_en & W0_addr_sel == 8'h6a;
  assign mem_106_3_W0_mask = W0_mask[3];
  assign mem_106_4_R0_addr = R0_addr[25:0];
  assign mem_106_4_R0_clk = R0_clk;
  assign mem_106_4_R0_en = R0_en & R0_addr_sel == 8'h6a;
  assign mem_106_4_W0_addr = W0_addr[25:0];
  assign mem_106_4_W0_clk = W0_clk;
  assign mem_106_4_W0_data = W0_data[39:32];
  assign mem_106_4_W0_en = W0_en & W0_addr_sel == 8'h6a;
  assign mem_106_4_W0_mask = W0_mask[4];
  assign mem_106_5_R0_addr = R0_addr[25:0];
  assign mem_106_5_R0_clk = R0_clk;
  assign mem_106_5_R0_en = R0_en & R0_addr_sel == 8'h6a;
  assign mem_106_5_W0_addr = W0_addr[25:0];
  assign mem_106_5_W0_clk = W0_clk;
  assign mem_106_5_W0_data = W0_data[47:40];
  assign mem_106_5_W0_en = W0_en & W0_addr_sel == 8'h6a;
  assign mem_106_5_W0_mask = W0_mask[5];
  assign mem_106_6_R0_addr = R0_addr[25:0];
  assign mem_106_6_R0_clk = R0_clk;
  assign mem_106_6_R0_en = R0_en & R0_addr_sel == 8'h6a;
  assign mem_106_6_W0_addr = W0_addr[25:0];
  assign mem_106_6_W0_clk = W0_clk;
  assign mem_106_6_W0_data = W0_data[55:48];
  assign mem_106_6_W0_en = W0_en & W0_addr_sel == 8'h6a;
  assign mem_106_6_W0_mask = W0_mask[6];
  assign mem_106_7_R0_addr = R0_addr[25:0];
  assign mem_106_7_R0_clk = R0_clk;
  assign mem_106_7_R0_en = R0_en & R0_addr_sel == 8'h6a;
  assign mem_106_7_W0_addr = W0_addr[25:0];
  assign mem_106_7_W0_clk = W0_clk;
  assign mem_106_7_W0_data = W0_data[63:56];
  assign mem_106_7_W0_en = W0_en & W0_addr_sel == 8'h6a;
  assign mem_106_7_W0_mask = W0_mask[7];
  assign mem_107_0_R0_addr = R0_addr[25:0];
  assign mem_107_0_R0_clk = R0_clk;
  assign mem_107_0_R0_en = R0_en & R0_addr_sel == 8'h6b;
  assign mem_107_0_W0_addr = W0_addr[25:0];
  assign mem_107_0_W0_clk = W0_clk;
  assign mem_107_0_W0_data = W0_data[7:0];
  assign mem_107_0_W0_en = W0_en & W0_addr_sel == 8'h6b;
  assign mem_107_0_W0_mask = W0_mask[0];
  assign mem_107_1_R0_addr = R0_addr[25:0];
  assign mem_107_1_R0_clk = R0_clk;
  assign mem_107_1_R0_en = R0_en & R0_addr_sel == 8'h6b;
  assign mem_107_1_W0_addr = W0_addr[25:0];
  assign mem_107_1_W0_clk = W0_clk;
  assign mem_107_1_W0_data = W0_data[15:8];
  assign mem_107_1_W0_en = W0_en & W0_addr_sel == 8'h6b;
  assign mem_107_1_W0_mask = W0_mask[1];
  assign mem_107_2_R0_addr = R0_addr[25:0];
  assign mem_107_2_R0_clk = R0_clk;
  assign mem_107_2_R0_en = R0_en & R0_addr_sel == 8'h6b;
  assign mem_107_2_W0_addr = W0_addr[25:0];
  assign mem_107_2_W0_clk = W0_clk;
  assign mem_107_2_W0_data = W0_data[23:16];
  assign mem_107_2_W0_en = W0_en & W0_addr_sel == 8'h6b;
  assign mem_107_2_W0_mask = W0_mask[2];
  assign mem_107_3_R0_addr = R0_addr[25:0];
  assign mem_107_3_R0_clk = R0_clk;
  assign mem_107_3_R0_en = R0_en & R0_addr_sel == 8'h6b;
  assign mem_107_3_W0_addr = W0_addr[25:0];
  assign mem_107_3_W0_clk = W0_clk;
  assign mem_107_3_W0_data = W0_data[31:24];
  assign mem_107_3_W0_en = W0_en & W0_addr_sel == 8'h6b;
  assign mem_107_3_W0_mask = W0_mask[3];
  assign mem_107_4_R0_addr = R0_addr[25:0];
  assign mem_107_4_R0_clk = R0_clk;
  assign mem_107_4_R0_en = R0_en & R0_addr_sel == 8'h6b;
  assign mem_107_4_W0_addr = W0_addr[25:0];
  assign mem_107_4_W0_clk = W0_clk;
  assign mem_107_4_W0_data = W0_data[39:32];
  assign mem_107_4_W0_en = W0_en & W0_addr_sel == 8'h6b;
  assign mem_107_4_W0_mask = W0_mask[4];
  assign mem_107_5_R0_addr = R0_addr[25:0];
  assign mem_107_5_R0_clk = R0_clk;
  assign mem_107_5_R0_en = R0_en & R0_addr_sel == 8'h6b;
  assign mem_107_5_W0_addr = W0_addr[25:0];
  assign mem_107_5_W0_clk = W0_clk;
  assign mem_107_5_W0_data = W0_data[47:40];
  assign mem_107_5_W0_en = W0_en & W0_addr_sel == 8'h6b;
  assign mem_107_5_W0_mask = W0_mask[5];
  assign mem_107_6_R0_addr = R0_addr[25:0];
  assign mem_107_6_R0_clk = R0_clk;
  assign mem_107_6_R0_en = R0_en & R0_addr_sel == 8'h6b;
  assign mem_107_6_W0_addr = W0_addr[25:0];
  assign mem_107_6_W0_clk = W0_clk;
  assign mem_107_6_W0_data = W0_data[55:48];
  assign mem_107_6_W0_en = W0_en & W0_addr_sel == 8'h6b;
  assign mem_107_6_W0_mask = W0_mask[6];
  assign mem_107_7_R0_addr = R0_addr[25:0];
  assign mem_107_7_R0_clk = R0_clk;
  assign mem_107_7_R0_en = R0_en & R0_addr_sel == 8'h6b;
  assign mem_107_7_W0_addr = W0_addr[25:0];
  assign mem_107_7_W0_clk = W0_clk;
  assign mem_107_7_W0_data = W0_data[63:56];
  assign mem_107_7_W0_en = W0_en & W0_addr_sel == 8'h6b;
  assign mem_107_7_W0_mask = W0_mask[7];
  assign mem_108_0_R0_addr = R0_addr[25:0];
  assign mem_108_0_R0_clk = R0_clk;
  assign mem_108_0_R0_en = R0_en & R0_addr_sel == 8'h6c;
  assign mem_108_0_W0_addr = W0_addr[25:0];
  assign mem_108_0_W0_clk = W0_clk;
  assign mem_108_0_W0_data = W0_data[7:0];
  assign mem_108_0_W0_en = W0_en & W0_addr_sel == 8'h6c;
  assign mem_108_0_W0_mask = W0_mask[0];
  assign mem_108_1_R0_addr = R0_addr[25:0];
  assign mem_108_1_R0_clk = R0_clk;
  assign mem_108_1_R0_en = R0_en & R0_addr_sel == 8'h6c;
  assign mem_108_1_W0_addr = W0_addr[25:0];
  assign mem_108_1_W0_clk = W0_clk;
  assign mem_108_1_W0_data = W0_data[15:8];
  assign mem_108_1_W0_en = W0_en & W0_addr_sel == 8'h6c;
  assign mem_108_1_W0_mask = W0_mask[1];
  assign mem_108_2_R0_addr = R0_addr[25:0];
  assign mem_108_2_R0_clk = R0_clk;
  assign mem_108_2_R0_en = R0_en & R0_addr_sel == 8'h6c;
  assign mem_108_2_W0_addr = W0_addr[25:0];
  assign mem_108_2_W0_clk = W0_clk;
  assign mem_108_2_W0_data = W0_data[23:16];
  assign mem_108_2_W0_en = W0_en & W0_addr_sel == 8'h6c;
  assign mem_108_2_W0_mask = W0_mask[2];
  assign mem_108_3_R0_addr = R0_addr[25:0];
  assign mem_108_3_R0_clk = R0_clk;
  assign mem_108_3_R0_en = R0_en & R0_addr_sel == 8'h6c;
  assign mem_108_3_W0_addr = W0_addr[25:0];
  assign mem_108_3_W0_clk = W0_clk;
  assign mem_108_3_W0_data = W0_data[31:24];
  assign mem_108_3_W0_en = W0_en & W0_addr_sel == 8'h6c;
  assign mem_108_3_W0_mask = W0_mask[3];
  assign mem_108_4_R0_addr = R0_addr[25:0];
  assign mem_108_4_R0_clk = R0_clk;
  assign mem_108_4_R0_en = R0_en & R0_addr_sel == 8'h6c;
  assign mem_108_4_W0_addr = W0_addr[25:0];
  assign mem_108_4_W0_clk = W0_clk;
  assign mem_108_4_W0_data = W0_data[39:32];
  assign mem_108_4_W0_en = W0_en & W0_addr_sel == 8'h6c;
  assign mem_108_4_W0_mask = W0_mask[4];
  assign mem_108_5_R0_addr = R0_addr[25:0];
  assign mem_108_5_R0_clk = R0_clk;
  assign mem_108_5_R0_en = R0_en & R0_addr_sel == 8'h6c;
  assign mem_108_5_W0_addr = W0_addr[25:0];
  assign mem_108_5_W0_clk = W0_clk;
  assign mem_108_5_W0_data = W0_data[47:40];
  assign mem_108_5_W0_en = W0_en & W0_addr_sel == 8'h6c;
  assign mem_108_5_W0_mask = W0_mask[5];
  assign mem_108_6_R0_addr = R0_addr[25:0];
  assign mem_108_6_R0_clk = R0_clk;
  assign mem_108_6_R0_en = R0_en & R0_addr_sel == 8'h6c;
  assign mem_108_6_W0_addr = W0_addr[25:0];
  assign mem_108_6_W0_clk = W0_clk;
  assign mem_108_6_W0_data = W0_data[55:48];
  assign mem_108_6_W0_en = W0_en & W0_addr_sel == 8'h6c;
  assign mem_108_6_W0_mask = W0_mask[6];
  assign mem_108_7_R0_addr = R0_addr[25:0];
  assign mem_108_7_R0_clk = R0_clk;
  assign mem_108_7_R0_en = R0_en & R0_addr_sel == 8'h6c;
  assign mem_108_7_W0_addr = W0_addr[25:0];
  assign mem_108_7_W0_clk = W0_clk;
  assign mem_108_7_W0_data = W0_data[63:56];
  assign mem_108_7_W0_en = W0_en & W0_addr_sel == 8'h6c;
  assign mem_108_7_W0_mask = W0_mask[7];
  assign mem_109_0_R0_addr = R0_addr[25:0];
  assign mem_109_0_R0_clk = R0_clk;
  assign mem_109_0_R0_en = R0_en & R0_addr_sel == 8'h6d;
  assign mem_109_0_W0_addr = W0_addr[25:0];
  assign mem_109_0_W0_clk = W0_clk;
  assign mem_109_0_W0_data = W0_data[7:0];
  assign mem_109_0_W0_en = W0_en & W0_addr_sel == 8'h6d;
  assign mem_109_0_W0_mask = W0_mask[0];
  assign mem_109_1_R0_addr = R0_addr[25:0];
  assign mem_109_1_R0_clk = R0_clk;
  assign mem_109_1_R0_en = R0_en & R0_addr_sel == 8'h6d;
  assign mem_109_1_W0_addr = W0_addr[25:0];
  assign mem_109_1_W0_clk = W0_clk;
  assign mem_109_1_W0_data = W0_data[15:8];
  assign mem_109_1_W0_en = W0_en & W0_addr_sel == 8'h6d;
  assign mem_109_1_W0_mask = W0_mask[1];
  assign mem_109_2_R0_addr = R0_addr[25:0];
  assign mem_109_2_R0_clk = R0_clk;
  assign mem_109_2_R0_en = R0_en & R0_addr_sel == 8'h6d;
  assign mem_109_2_W0_addr = W0_addr[25:0];
  assign mem_109_2_W0_clk = W0_clk;
  assign mem_109_2_W0_data = W0_data[23:16];
  assign mem_109_2_W0_en = W0_en & W0_addr_sel == 8'h6d;
  assign mem_109_2_W0_mask = W0_mask[2];
  assign mem_109_3_R0_addr = R0_addr[25:0];
  assign mem_109_3_R0_clk = R0_clk;
  assign mem_109_3_R0_en = R0_en & R0_addr_sel == 8'h6d;
  assign mem_109_3_W0_addr = W0_addr[25:0];
  assign mem_109_3_W0_clk = W0_clk;
  assign mem_109_3_W0_data = W0_data[31:24];
  assign mem_109_3_W0_en = W0_en & W0_addr_sel == 8'h6d;
  assign mem_109_3_W0_mask = W0_mask[3];
  assign mem_109_4_R0_addr = R0_addr[25:0];
  assign mem_109_4_R0_clk = R0_clk;
  assign mem_109_4_R0_en = R0_en & R0_addr_sel == 8'h6d;
  assign mem_109_4_W0_addr = W0_addr[25:0];
  assign mem_109_4_W0_clk = W0_clk;
  assign mem_109_4_W0_data = W0_data[39:32];
  assign mem_109_4_W0_en = W0_en & W0_addr_sel == 8'h6d;
  assign mem_109_4_W0_mask = W0_mask[4];
  assign mem_109_5_R0_addr = R0_addr[25:0];
  assign mem_109_5_R0_clk = R0_clk;
  assign mem_109_5_R0_en = R0_en & R0_addr_sel == 8'h6d;
  assign mem_109_5_W0_addr = W0_addr[25:0];
  assign mem_109_5_W0_clk = W0_clk;
  assign mem_109_5_W0_data = W0_data[47:40];
  assign mem_109_5_W0_en = W0_en & W0_addr_sel == 8'h6d;
  assign mem_109_5_W0_mask = W0_mask[5];
  assign mem_109_6_R0_addr = R0_addr[25:0];
  assign mem_109_6_R0_clk = R0_clk;
  assign mem_109_6_R0_en = R0_en & R0_addr_sel == 8'h6d;
  assign mem_109_6_W0_addr = W0_addr[25:0];
  assign mem_109_6_W0_clk = W0_clk;
  assign mem_109_6_W0_data = W0_data[55:48];
  assign mem_109_6_W0_en = W0_en & W0_addr_sel == 8'h6d;
  assign mem_109_6_W0_mask = W0_mask[6];
  assign mem_109_7_R0_addr = R0_addr[25:0];
  assign mem_109_7_R0_clk = R0_clk;
  assign mem_109_7_R0_en = R0_en & R0_addr_sel == 8'h6d;
  assign mem_109_7_W0_addr = W0_addr[25:0];
  assign mem_109_7_W0_clk = W0_clk;
  assign mem_109_7_W0_data = W0_data[63:56];
  assign mem_109_7_W0_en = W0_en & W0_addr_sel == 8'h6d;
  assign mem_109_7_W0_mask = W0_mask[7];
  assign mem_110_0_R0_addr = R0_addr[25:0];
  assign mem_110_0_R0_clk = R0_clk;
  assign mem_110_0_R0_en = R0_en & R0_addr_sel == 8'h6e;
  assign mem_110_0_W0_addr = W0_addr[25:0];
  assign mem_110_0_W0_clk = W0_clk;
  assign mem_110_0_W0_data = W0_data[7:0];
  assign mem_110_0_W0_en = W0_en & W0_addr_sel == 8'h6e;
  assign mem_110_0_W0_mask = W0_mask[0];
  assign mem_110_1_R0_addr = R0_addr[25:0];
  assign mem_110_1_R0_clk = R0_clk;
  assign mem_110_1_R0_en = R0_en & R0_addr_sel == 8'h6e;
  assign mem_110_1_W0_addr = W0_addr[25:0];
  assign mem_110_1_W0_clk = W0_clk;
  assign mem_110_1_W0_data = W0_data[15:8];
  assign mem_110_1_W0_en = W0_en & W0_addr_sel == 8'h6e;
  assign mem_110_1_W0_mask = W0_mask[1];
  assign mem_110_2_R0_addr = R0_addr[25:0];
  assign mem_110_2_R0_clk = R0_clk;
  assign mem_110_2_R0_en = R0_en & R0_addr_sel == 8'h6e;
  assign mem_110_2_W0_addr = W0_addr[25:0];
  assign mem_110_2_W0_clk = W0_clk;
  assign mem_110_2_W0_data = W0_data[23:16];
  assign mem_110_2_W0_en = W0_en & W0_addr_sel == 8'h6e;
  assign mem_110_2_W0_mask = W0_mask[2];
  assign mem_110_3_R0_addr = R0_addr[25:0];
  assign mem_110_3_R0_clk = R0_clk;
  assign mem_110_3_R0_en = R0_en & R0_addr_sel == 8'h6e;
  assign mem_110_3_W0_addr = W0_addr[25:0];
  assign mem_110_3_W0_clk = W0_clk;
  assign mem_110_3_W0_data = W0_data[31:24];
  assign mem_110_3_W0_en = W0_en & W0_addr_sel == 8'h6e;
  assign mem_110_3_W0_mask = W0_mask[3];
  assign mem_110_4_R0_addr = R0_addr[25:0];
  assign mem_110_4_R0_clk = R0_clk;
  assign mem_110_4_R0_en = R0_en & R0_addr_sel == 8'h6e;
  assign mem_110_4_W0_addr = W0_addr[25:0];
  assign mem_110_4_W0_clk = W0_clk;
  assign mem_110_4_W0_data = W0_data[39:32];
  assign mem_110_4_W0_en = W0_en & W0_addr_sel == 8'h6e;
  assign mem_110_4_W0_mask = W0_mask[4];
  assign mem_110_5_R0_addr = R0_addr[25:0];
  assign mem_110_5_R0_clk = R0_clk;
  assign mem_110_5_R0_en = R0_en & R0_addr_sel == 8'h6e;
  assign mem_110_5_W0_addr = W0_addr[25:0];
  assign mem_110_5_W0_clk = W0_clk;
  assign mem_110_5_W0_data = W0_data[47:40];
  assign mem_110_5_W0_en = W0_en & W0_addr_sel == 8'h6e;
  assign mem_110_5_W0_mask = W0_mask[5];
  assign mem_110_6_R0_addr = R0_addr[25:0];
  assign mem_110_6_R0_clk = R0_clk;
  assign mem_110_6_R0_en = R0_en & R0_addr_sel == 8'h6e;
  assign mem_110_6_W0_addr = W0_addr[25:0];
  assign mem_110_6_W0_clk = W0_clk;
  assign mem_110_6_W0_data = W0_data[55:48];
  assign mem_110_6_W0_en = W0_en & W0_addr_sel == 8'h6e;
  assign mem_110_6_W0_mask = W0_mask[6];
  assign mem_110_7_R0_addr = R0_addr[25:0];
  assign mem_110_7_R0_clk = R0_clk;
  assign mem_110_7_R0_en = R0_en & R0_addr_sel == 8'h6e;
  assign mem_110_7_W0_addr = W0_addr[25:0];
  assign mem_110_7_W0_clk = W0_clk;
  assign mem_110_7_W0_data = W0_data[63:56];
  assign mem_110_7_W0_en = W0_en & W0_addr_sel == 8'h6e;
  assign mem_110_7_W0_mask = W0_mask[7];
  assign mem_111_0_R0_addr = R0_addr[25:0];
  assign mem_111_0_R0_clk = R0_clk;
  assign mem_111_0_R0_en = R0_en & R0_addr_sel == 8'h6f;
  assign mem_111_0_W0_addr = W0_addr[25:0];
  assign mem_111_0_W0_clk = W0_clk;
  assign mem_111_0_W0_data = W0_data[7:0];
  assign mem_111_0_W0_en = W0_en & W0_addr_sel == 8'h6f;
  assign mem_111_0_W0_mask = W0_mask[0];
  assign mem_111_1_R0_addr = R0_addr[25:0];
  assign mem_111_1_R0_clk = R0_clk;
  assign mem_111_1_R0_en = R0_en & R0_addr_sel == 8'h6f;
  assign mem_111_1_W0_addr = W0_addr[25:0];
  assign mem_111_1_W0_clk = W0_clk;
  assign mem_111_1_W0_data = W0_data[15:8];
  assign mem_111_1_W0_en = W0_en & W0_addr_sel == 8'h6f;
  assign mem_111_1_W0_mask = W0_mask[1];
  assign mem_111_2_R0_addr = R0_addr[25:0];
  assign mem_111_2_R0_clk = R0_clk;
  assign mem_111_2_R0_en = R0_en & R0_addr_sel == 8'h6f;
  assign mem_111_2_W0_addr = W0_addr[25:0];
  assign mem_111_2_W0_clk = W0_clk;
  assign mem_111_2_W0_data = W0_data[23:16];
  assign mem_111_2_W0_en = W0_en & W0_addr_sel == 8'h6f;
  assign mem_111_2_W0_mask = W0_mask[2];
  assign mem_111_3_R0_addr = R0_addr[25:0];
  assign mem_111_3_R0_clk = R0_clk;
  assign mem_111_3_R0_en = R0_en & R0_addr_sel == 8'h6f;
  assign mem_111_3_W0_addr = W0_addr[25:0];
  assign mem_111_3_W0_clk = W0_clk;
  assign mem_111_3_W0_data = W0_data[31:24];
  assign mem_111_3_W0_en = W0_en & W0_addr_sel == 8'h6f;
  assign mem_111_3_W0_mask = W0_mask[3];
  assign mem_111_4_R0_addr = R0_addr[25:0];
  assign mem_111_4_R0_clk = R0_clk;
  assign mem_111_4_R0_en = R0_en & R0_addr_sel == 8'h6f;
  assign mem_111_4_W0_addr = W0_addr[25:0];
  assign mem_111_4_W0_clk = W0_clk;
  assign mem_111_4_W0_data = W0_data[39:32];
  assign mem_111_4_W0_en = W0_en & W0_addr_sel == 8'h6f;
  assign mem_111_4_W0_mask = W0_mask[4];
  assign mem_111_5_R0_addr = R0_addr[25:0];
  assign mem_111_5_R0_clk = R0_clk;
  assign mem_111_5_R0_en = R0_en & R0_addr_sel == 8'h6f;
  assign mem_111_5_W0_addr = W0_addr[25:0];
  assign mem_111_5_W0_clk = W0_clk;
  assign mem_111_5_W0_data = W0_data[47:40];
  assign mem_111_5_W0_en = W0_en & W0_addr_sel == 8'h6f;
  assign mem_111_5_W0_mask = W0_mask[5];
  assign mem_111_6_R0_addr = R0_addr[25:0];
  assign mem_111_6_R0_clk = R0_clk;
  assign mem_111_6_R0_en = R0_en & R0_addr_sel == 8'h6f;
  assign mem_111_6_W0_addr = W0_addr[25:0];
  assign mem_111_6_W0_clk = W0_clk;
  assign mem_111_6_W0_data = W0_data[55:48];
  assign mem_111_6_W0_en = W0_en & W0_addr_sel == 8'h6f;
  assign mem_111_6_W0_mask = W0_mask[6];
  assign mem_111_7_R0_addr = R0_addr[25:0];
  assign mem_111_7_R0_clk = R0_clk;
  assign mem_111_7_R0_en = R0_en & R0_addr_sel == 8'h6f;
  assign mem_111_7_W0_addr = W0_addr[25:0];
  assign mem_111_7_W0_clk = W0_clk;
  assign mem_111_7_W0_data = W0_data[63:56];
  assign mem_111_7_W0_en = W0_en & W0_addr_sel == 8'h6f;
  assign mem_111_7_W0_mask = W0_mask[7];
  assign mem_112_0_R0_addr = R0_addr[25:0];
  assign mem_112_0_R0_clk = R0_clk;
  assign mem_112_0_R0_en = R0_en & R0_addr_sel == 8'h70;
  assign mem_112_0_W0_addr = W0_addr[25:0];
  assign mem_112_0_W0_clk = W0_clk;
  assign mem_112_0_W0_data = W0_data[7:0];
  assign mem_112_0_W0_en = W0_en & W0_addr_sel == 8'h70;
  assign mem_112_0_W0_mask = W0_mask[0];
  assign mem_112_1_R0_addr = R0_addr[25:0];
  assign mem_112_1_R0_clk = R0_clk;
  assign mem_112_1_R0_en = R0_en & R0_addr_sel == 8'h70;
  assign mem_112_1_W0_addr = W0_addr[25:0];
  assign mem_112_1_W0_clk = W0_clk;
  assign mem_112_1_W0_data = W0_data[15:8];
  assign mem_112_1_W0_en = W0_en & W0_addr_sel == 8'h70;
  assign mem_112_1_W0_mask = W0_mask[1];
  assign mem_112_2_R0_addr = R0_addr[25:0];
  assign mem_112_2_R0_clk = R0_clk;
  assign mem_112_2_R0_en = R0_en & R0_addr_sel == 8'h70;
  assign mem_112_2_W0_addr = W0_addr[25:0];
  assign mem_112_2_W0_clk = W0_clk;
  assign mem_112_2_W0_data = W0_data[23:16];
  assign mem_112_2_W0_en = W0_en & W0_addr_sel == 8'h70;
  assign mem_112_2_W0_mask = W0_mask[2];
  assign mem_112_3_R0_addr = R0_addr[25:0];
  assign mem_112_3_R0_clk = R0_clk;
  assign mem_112_3_R0_en = R0_en & R0_addr_sel == 8'h70;
  assign mem_112_3_W0_addr = W0_addr[25:0];
  assign mem_112_3_W0_clk = W0_clk;
  assign mem_112_3_W0_data = W0_data[31:24];
  assign mem_112_3_W0_en = W0_en & W0_addr_sel == 8'h70;
  assign mem_112_3_W0_mask = W0_mask[3];
  assign mem_112_4_R0_addr = R0_addr[25:0];
  assign mem_112_4_R0_clk = R0_clk;
  assign mem_112_4_R0_en = R0_en & R0_addr_sel == 8'h70;
  assign mem_112_4_W0_addr = W0_addr[25:0];
  assign mem_112_4_W0_clk = W0_clk;
  assign mem_112_4_W0_data = W0_data[39:32];
  assign mem_112_4_W0_en = W0_en & W0_addr_sel == 8'h70;
  assign mem_112_4_W0_mask = W0_mask[4];
  assign mem_112_5_R0_addr = R0_addr[25:0];
  assign mem_112_5_R0_clk = R0_clk;
  assign mem_112_5_R0_en = R0_en & R0_addr_sel == 8'h70;
  assign mem_112_5_W0_addr = W0_addr[25:0];
  assign mem_112_5_W0_clk = W0_clk;
  assign mem_112_5_W0_data = W0_data[47:40];
  assign mem_112_5_W0_en = W0_en & W0_addr_sel == 8'h70;
  assign mem_112_5_W0_mask = W0_mask[5];
  assign mem_112_6_R0_addr = R0_addr[25:0];
  assign mem_112_6_R0_clk = R0_clk;
  assign mem_112_6_R0_en = R0_en & R0_addr_sel == 8'h70;
  assign mem_112_6_W0_addr = W0_addr[25:0];
  assign mem_112_6_W0_clk = W0_clk;
  assign mem_112_6_W0_data = W0_data[55:48];
  assign mem_112_6_W0_en = W0_en & W0_addr_sel == 8'h70;
  assign mem_112_6_W0_mask = W0_mask[6];
  assign mem_112_7_R0_addr = R0_addr[25:0];
  assign mem_112_7_R0_clk = R0_clk;
  assign mem_112_7_R0_en = R0_en & R0_addr_sel == 8'h70;
  assign mem_112_7_W0_addr = W0_addr[25:0];
  assign mem_112_7_W0_clk = W0_clk;
  assign mem_112_7_W0_data = W0_data[63:56];
  assign mem_112_7_W0_en = W0_en & W0_addr_sel == 8'h70;
  assign mem_112_7_W0_mask = W0_mask[7];
  assign mem_113_0_R0_addr = R0_addr[25:0];
  assign mem_113_0_R0_clk = R0_clk;
  assign mem_113_0_R0_en = R0_en & R0_addr_sel == 8'h71;
  assign mem_113_0_W0_addr = W0_addr[25:0];
  assign mem_113_0_W0_clk = W0_clk;
  assign mem_113_0_W0_data = W0_data[7:0];
  assign mem_113_0_W0_en = W0_en & W0_addr_sel == 8'h71;
  assign mem_113_0_W0_mask = W0_mask[0];
  assign mem_113_1_R0_addr = R0_addr[25:0];
  assign mem_113_1_R0_clk = R0_clk;
  assign mem_113_1_R0_en = R0_en & R0_addr_sel == 8'h71;
  assign mem_113_1_W0_addr = W0_addr[25:0];
  assign mem_113_1_W0_clk = W0_clk;
  assign mem_113_1_W0_data = W0_data[15:8];
  assign mem_113_1_W0_en = W0_en & W0_addr_sel == 8'h71;
  assign mem_113_1_W0_mask = W0_mask[1];
  assign mem_113_2_R0_addr = R0_addr[25:0];
  assign mem_113_2_R0_clk = R0_clk;
  assign mem_113_2_R0_en = R0_en & R0_addr_sel == 8'h71;
  assign mem_113_2_W0_addr = W0_addr[25:0];
  assign mem_113_2_W0_clk = W0_clk;
  assign mem_113_2_W0_data = W0_data[23:16];
  assign mem_113_2_W0_en = W0_en & W0_addr_sel == 8'h71;
  assign mem_113_2_W0_mask = W0_mask[2];
  assign mem_113_3_R0_addr = R0_addr[25:0];
  assign mem_113_3_R0_clk = R0_clk;
  assign mem_113_3_R0_en = R0_en & R0_addr_sel == 8'h71;
  assign mem_113_3_W0_addr = W0_addr[25:0];
  assign mem_113_3_W0_clk = W0_clk;
  assign mem_113_3_W0_data = W0_data[31:24];
  assign mem_113_3_W0_en = W0_en & W0_addr_sel == 8'h71;
  assign mem_113_3_W0_mask = W0_mask[3];
  assign mem_113_4_R0_addr = R0_addr[25:0];
  assign mem_113_4_R0_clk = R0_clk;
  assign mem_113_4_R0_en = R0_en & R0_addr_sel == 8'h71;
  assign mem_113_4_W0_addr = W0_addr[25:0];
  assign mem_113_4_W0_clk = W0_clk;
  assign mem_113_4_W0_data = W0_data[39:32];
  assign mem_113_4_W0_en = W0_en & W0_addr_sel == 8'h71;
  assign mem_113_4_W0_mask = W0_mask[4];
  assign mem_113_5_R0_addr = R0_addr[25:0];
  assign mem_113_5_R0_clk = R0_clk;
  assign mem_113_5_R0_en = R0_en & R0_addr_sel == 8'h71;
  assign mem_113_5_W0_addr = W0_addr[25:0];
  assign mem_113_5_W0_clk = W0_clk;
  assign mem_113_5_W0_data = W0_data[47:40];
  assign mem_113_5_W0_en = W0_en & W0_addr_sel == 8'h71;
  assign mem_113_5_W0_mask = W0_mask[5];
  assign mem_113_6_R0_addr = R0_addr[25:0];
  assign mem_113_6_R0_clk = R0_clk;
  assign mem_113_6_R0_en = R0_en & R0_addr_sel == 8'h71;
  assign mem_113_6_W0_addr = W0_addr[25:0];
  assign mem_113_6_W0_clk = W0_clk;
  assign mem_113_6_W0_data = W0_data[55:48];
  assign mem_113_6_W0_en = W0_en & W0_addr_sel == 8'h71;
  assign mem_113_6_W0_mask = W0_mask[6];
  assign mem_113_7_R0_addr = R0_addr[25:0];
  assign mem_113_7_R0_clk = R0_clk;
  assign mem_113_7_R0_en = R0_en & R0_addr_sel == 8'h71;
  assign mem_113_7_W0_addr = W0_addr[25:0];
  assign mem_113_7_W0_clk = W0_clk;
  assign mem_113_7_W0_data = W0_data[63:56];
  assign mem_113_7_W0_en = W0_en & W0_addr_sel == 8'h71;
  assign mem_113_7_W0_mask = W0_mask[7];
  assign mem_114_0_R0_addr = R0_addr[25:0];
  assign mem_114_0_R0_clk = R0_clk;
  assign mem_114_0_R0_en = R0_en & R0_addr_sel == 8'h72;
  assign mem_114_0_W0_addr = W0_addr[25:0];
  assign mem_114_0_W0_clk = W0_clk;
  assign mem_114_0_W0_data = W0_data[7:0];
  assign mem_114_0_W0_en = W0_en & W0_addr_sel == 8'h72;
  assign mem_114_0_W0_mask = W0_mask[0];
  assign mem_114_1_R0_addr = R0_addr[25:0];
  assign mem_114_1_R0_clk = R0_clk;
  assign mem_114_1_R0_en = R0_en & R0_addr_sel == 8'h72;
  assign mem_114_1_W0_addr = W0_addr[25:0];
  assign mem_114_1_W0_clk = W0_clk;
  assign mem_114_1_W0_data = W0_data[15:8];
  assign mem_114_1_W0_en = W0_en & W0_addr_sel == 8'h72;
  assign mem_114_1_W0_mask = W0_mask[1];
  assign mem_114_2_R0_addr = R0_addr[25:0];
  assign mem_114_2_R0_clk = R0_clk;
  assign mem_114_2_R0_en = R0_en & R0_addr_sel == 8'h72;
  assign mem_114_2_W0_addr = W0_addr[25:0];
  assign mem_114_2_W0_clk = W0_clk;
  assign mem_114_2_W0_data = W0_data[23:16];
  assign mem_114_2_W0_en = W0_en & W0_addr_sel == 8'h72;
  assign mem_114_2_W0_mask = W0_mask[2];
  assign mem_114_3_R0_addr = R0_addr[25:0];
  assign mem_114_3_R0_clk = R0_clk;
  assign mem_114_3_R0_en = R0_en & R0_addr_sel == 8'h72;
  assign mem_114_3_W0_addr = W0_addr[25:0];
  assign mem_114_3_W0_clk = W0_clk;
  assign mem_114_3_W0_data = W0_data[31:24];
  assign mem_114_3_W0_en = W0_en & W0_addr_sel == 8'h72;
  assign mem_114_3_W0_mask = W0_mask[3];
  assign mem_114_4_R0_addr = R0_addr[25:0];
  assign mem_114_4_R0_clk = R0_clk;
  assign mem_114_4_R0_en = R0_en & R0_addr_sel == 8'h72;
  assign mem_114_4_W0_addr = W0_addr[25:0];
  assign mem_114_4_W0_clk = W0_clk;
  assign mem_114_4_W0_data = W0_data[39:32];
  assign mem_114_4_W0_en = W0_en & W0_addr_sel == 8'h72;
  assign mem_114_4_W0_mask = W0_mask[4];
  assign mem_114_5_R0_addr = R0_addr[25:0];
  assign mem_114_5_R0_clk = R0_clk;
  assign mem_114_5_R0_en = R0_en & R0_addr_sel == 8'h72;
  assign mem_114_5_W0_addr = W0_addr[25:0];
  assign mem_114_5_W0_clk = W0_clk;
  assign mem_114_5_W0_data = W0_data[47:40];
  assign mem_114_5_W0_en = W0_en & W0_addr_sel == 8'h72;
  assign mem_114_5_W0_mask = W0_mask[5];
  assign mem_114_6_R0_addr = R0_addr[25:0];
  assign mem_114_6_R0_clk = R0_clk;
  assign mem_114_6_R0_en = R0_en & R0_addr_sel == 8'h72;
  assign mem_114_6_W0_addr = W0_addr[25:0];
  assign mem_114_6_W0_clk = W0_clk;
  assign mem_114_6_W0_data = W0_data[55:48];
  assign mem_114_6_W0_en = W0_en & W0_addr_sel == 8'h72;
  assign mem_114_6_W0_mask = W0_mask[6];
  assign mem_114_7_R0_addr = R0_addr[25:0];
  assign mem_114_7_R0_clk = R0_clk;
  assign mem_114_7_R0_en = R0_en & R0_addr_sel == 8'h72;
  assign mem_114_7_W0_addr = W0_addr[25:0];
  assign mem_114_7_W0_clk = W0_clk;
  assign mem_114_7_W0_data = W0_data[63:56];
  assign mem_114_7_W0_en = W0_en & W0_addr_sel == 8'h72;
  assign mem_114_7_W0_mask = W0_mask[7];
  assign mem_115_0_R0_addr = R0_addr[25:0];
  assign mem_115_0_R0_clk = R0_clk;
  assign mem_115_0_R0_en = R0_en & R0_addr_sel == 8'h73;
  assign mem_115_0_W0_addr = W0_addr[25:0];
  assign mem_115_0_W0_clk = W0_clk;
  assign mem_115_0_W0_data = W0_data[7:0];
  assign mem_115_0_W0_en = W0_en & W0_addr_sel == 8'h73;
  assign mem_115_0_W0_mask = W0_mask[0];
  assign mem_115_1_R0_addr = R0_addr[25:0];
  assign mem_115_1_R0_clk = R0_clk;
  assign mem_115_1_R0_en = R0_en & R0_addr_sel == 8'h73;
  assign mem_115_1_W0_addr = W0_addr[25:0];
  assign mem_115_1_W0_clk = W0_clk;
  assign mem_115_1_W0_data = W0_data[15:8];
  assign mem_115_1_W0_en = W0_en & W0_addr_sel == 8'h73;
  assign mem_115_1_W0_mask = W0_mask[1];
  assign mem_115_2_R0_addr = R0_addr[25:0];
  assign mem_115_2_R0_clk = R0_clk;
  assign mem_115_2_R0_en = R0_en & R0_addr_sel == 8'h73;
  assign mem_115_2_W0_addr = W0_addr[25:0];
  assign mem_115_2_W0_clk = W0_clk;
  assign mem_115_2_W0_data = W0_data[23:16];
  assign mem_115_2_W0_en = W0_en & W0_addr_sel == 8'h73;
  assign mem_115_2_W0_mask = W0_mask[2];
  assign mem_115_3_R0_addr = R0_addr[25:0];
  assign mem_115_3_R0_clk = R0_clk;
  assign mem_115_3_R0_en = R0_en & R0_addr_sel == 8'h73;
  assign mem_115_3_W0_addr = W0_addr[25:0];
  assign mem_115_3_W0_clk = W0_clk;
  assign mem_115_3_W0_data = W0_data[31:24];
  assign mem_115_3_W0_en = W0_en & W0_addr_sel == 8'h73;
  assign mem_115_3_W0_mask = W0_mask[3];
  assign mem_115_4_R0_addr = R0_addr[25:0];
  assign mem_115_4_R0_clk = R0_clk;
  assign mem_115_4_R0_en = R0_en & R0_addr_sel == 8'h73;
  assign mem_115_4_W0_addr = W0_addr[25:0];
  assign mem_115_4_W0_clk = W0_clk;
  assign mem_115_4_W0_data = W0_data[39:32];
  assign mem_115_4_W0_en = W0_en & W0_addr_sel == 8'h73;
  assign mem_115_4_W0_mask = W0_mask[4];
  assign mem_115_5_R0_addr = R0_addr[25:0];
  assign mem_115_5_R0_clk = R0_clk;
  assign mem_115_5_R0_en = R0_en & R0_addr_sel == 8'h73;
  assign mem_115_5_W0_addr = W0_addr[25:0];
  assign mem_115_5_W0_clk = W0_clk;
  assign mem_115_5_W0_data = W0_data[47:40];
  assign mem_115_5_W0_en = W0_en & W0_addr_sel == 8'h73;
  assign mem_115_5_W0_mask = W0_mask[5];
  assign mem_115_6_R0_addr = R0_addr[25:0];
  assign mem_115_6_R0_clk = R0_clk;
  assign mem_115_6_R0_en = R0_en & R0_addr_sel == 8'h73;
  assign mem_115_6_W0_addr = W0_addr[25:0];
  assign mem_115_6_W0_clk = W0_clk;
  assign mem_115_6_W0_data = W0_data[55:48];
  assign mem_115_6_W0_en = W0_en & W0_addr_sel == 8'h73;
  assign mem_115_6_W0_mask = W0_mask[6];
  assign mem_115_7_R0_addr = R0_addr[25:0];
  assign mem_115_7_R0_clk = R0_clk;
  assign mem_115_7_R0_en = R0_en & R0_addr_sel == 8'h73;
  assign mem_115_7_W0_addr = W0_addr[25:0];
  assign mem_115_7_W0_clk = W0_clk;
  assign mem_115_7_W0_data = W0_data[63:56];
  assign mem_115_7_W0_en = W0_en & W0_addr_sel == 8'h73;
  assign mem_115_7_W0_mask = W0_mask[7];
  assign mem_116_0_R0_addr = R0_addr[25:0];
  assign mem_116_0_R0_clk = R0_clk;
  assign mem_116_0_R0_en = R0_en & R0_addr_sel == 8'h74;
  assign mem_116_0_W0_addr = W0_addr[25:0];
  assign mem_116_0_W0_clk = W0_clk;
  assign mem_116_0_W0_data = W0_data[7:0];
  assign mem_116_0_W0_en = W0_en & W0_addr_sel == 8'h74;
  assign mem_116_0_W0_mask = W0_mask[0];
  assign mem_116_1_R0_addr = R0_addr[25:0];
  assign mem_116_1_R0_clk = R0_clk;
  assign mem_116_1_R0_en = R0_en & R0_addr_sel == 8'h74;
  assign mem_116_1_W0_addr = W0_addr[25:0];
  assign mem_116_1_W0_clk = W0_clk;
  assign mem_116_1_W0_data = W0_data[15:8];
  assign mem_116_1_W0_en = W0_en & W0_addr_sel == 8'h74;
  assign mem_116_1_W0_mask = W0_mask[1];
  assign mem_116_2_R0_addr = R0_addr[25:0];
  assign mem_116_2_R0_clk = R0_clk;
  assign mem_116_2_R0_en = R0_en & R0_addr_sel == 8'h74;
  assign mem_116_2_W0_addr = W0_addr[25:0];
  assign mem_116_2_W0_clk = W0_clk;
  assign mem_116_2_W0_data = W0_data[23:16];
  assign mem_116_2_W0_en = W0_en & W0_addr_sel == 8'h74;
  assign mem_116_2_W0_mask = W0_mask[2];
  assign mem_116_3_R0_addr = R0_addr[25:0];
  assign mem_116_3_R0_clk = R0_clk;
  assign mem_116_3_R0_en = R0_en & R0_addr_sel == 8'h74;
  assign mem_116_3_W0_addr = W0_addr[25:0];
  assign mem_116_3_W0_clk = W0_clk;
  assign mem_116_3_W0_data = W0_data[31:24];
  assign mem_116_3_W0_en = W0_en & W0_addr_sel == 8'h74;
  assign mem_116_3_W0_mask = W0_mask[3];
  assign mem_116_4_R0_addr = R0_addr[25:0];
  assign mem_116_4_R0_clk = R0_clk;
  assign mem_116_4_R0_en = R0_en & R0_addr_sel == 8'h74;
  assign mem_116_4_W0_addr = W0_addr[25:0];
  assign mem_116_4_W0_clk = W0_clk;
  assign mem_116_4_W0_data = W0_data[39:32];
  assign mem_116_4_W0_en = W0_en & W0_addr_sel == 8'h74;
  assign mem_116_4_W0_mask = W0_mask[4];
  assign mem_116_5_R0_addr = R0_addr[25:0];
  assign mem_116_5_R0_clk = R0_clk;
  assign mem_116_5_R0_en = R0_en & R0_addr_sel == 8'h74;
  assign mem_116_5_W0_addr = W0_addr[25:0];
  assign mem_116_5_W0_clk = W0_clk;
  assign mem_116_5_W0_data = W0_data[47:40];
  assign mem_116_5_W0_en = W0_en & W0_addr_sel == 8'h74;
  assign mem_116_5_W0_mask = W0_mask[5];
  assign mem_116_6_R0_addr = R0_addr[25:0];
  assign mem_116_6_R0_clk = R0_clk;
  assign mem_116_6_R0_en = R0_en & R0_addr_sel == 8'h74;
  assign mem_116_6_W0_addr = W0_addr[25:0];
  assign mem_116_6_W0_clk = W0_clk;
  assign mem_116_6_W0_data = W0_data[55:48];
  assign mem_116_6_W0_en = W0_en & W0_addr_sel == 8'h74;
  assign mem_116_6_W0_mask = W0_mask[6];
  assign mem_116_7_R0_addr = R0_addr[25:0];
  assign mem_116_7_R0_clk = R0_clk;
  assign mem_116_7_R0_en = R0_en & R0_addr_sel == 8'h74;
  assign mem_116_7_W0_addr = W0_addr[25:0];
  assign mem_116_7_W0_clk = W0_clk;
  assign mem_116_7_W0_data = W0_data[63:56];
  assign mem_116_7_W0_en = W0_en & W0_addr_sel == 8'h74;
  assign mem_116_7_W0_mask = W0_mask[7];
  assign mem_117_0_R0_addr = R0_addr[25:0];
  assign mem_117_0_R0_clk = R0_clk;
  assign mem_117_0_R0_en = R0_en & R0_addr_sel == 8'h75;
  assign mem_117_0_W0_addr = W0_addr[25:0];
  assign mem_117_0_W0_clk = W0_clk;
  assign mem_117_0_W0_data = W0_data[7:0];
  assign mem_117_0_W0_en = W0_en & W0_addr_sel == 8'h75;
  assign mem_117_0_W0_mask = W0_mask[0];
  assign mem_117_1_R0_addr = R0_addr[25:0];
  assign mem_117_1_R0_clk = R0_clk;
  assign mem_117_1_R0_en = R0_en & R0_addr_sel == 8'h75;
  assign mem_117_1_W0_addr = W0_addr[25:0];
  assign mem_117_1_W0_clk = W0_clk;
  assign mem_117_1_W0_data = W0_data[15:8];
  assign mem_117_1_W0_en = W0_en & W0_addr_sel == 8'h75;
  assign mem_117_1_W0_mask = W0_mask[1];
  assign mem_117_2_R0_addr = R0_addr[25:0];
  assign mem_117_2_R0_clk = R0_clk;
  assign mem_117_2_R0_en = R0_en & R0_addr_sel == 8'h75;
  assign mem_117_2_W0_addr = W0_addr[25:0];
  assign mem_117_2_W0_clk = W0_clk;
  assign mem_117_2_W0_data = W0_data[23:16];
  assign mem_117_2_W0_en = W0_en & W0_addr_sel == 8'h75;
  assign mem_117_2_W0_mask = W0_mask[2];
  assign mem_117_3_R0_addr = R0_addr[25:0];
  assign mem_117_3_R0_clk = R0_clk;
  assign mem_117_3_R0_en = R0_en & R0_addr_sel == 8'h75;
  assign mem_117_3_W0_addr = W0_addr[25:0];
  assign mem_117_3_W0_clk = W0_clk;
  assign mem_117_3_W0_data = W0_data[31:24];
  assign mem_117_3_W0_en = W0_en & W0_addr_sel == 8'h75;
  assign mem_117_3_W0_mask = W0_mask[3];
  assign mem_117_4_R0_addr = R0_addr[25:0];
  assign mem_117_4_R0_clk = R0_clk;
  assign mem_117_4_R0_en = R0_en & R0_addr_sel == 8'h75;
  assign mem_117_4_W0_addr = W0_addr[25:0];
  assign mem_117_4_W0_clk = W0_clk;
  assign mem_117_4_W0_data = W0_data[39:32];
  assign mem_117_4_W0_en = W0_en & W0_addr_sel == 8'h75;
  assign mem_117_4_W0_mask = W0_mask[4];
  assign mem_117_5_R0_addr = R0_addr[25:0];
  assign mem_117_5_R0_clk = R0_clk;
  assign mem_117_5_R0_en = R0_en & R0_addr_sel == 8'h75;
  assign mem_117_5_W0_addr = W0_addr[25:0];
  assign mem_117_5_W0_clk = W0_clk;
  assign mem_117_5_W0_data = W0_data[47:40];
  assign mem_117_5_W0_en = W0_en & W0_addr_sel == 8'h75;
  assign mem_117_5_W0_mask = W0_mask[5];
  assign mem_117_6_R0_addr = R0_addr[25:0];
  assign mem_117_6_R0_clk = R0_clk;
  assign mem_117_6_R0_en = R0_en & R0_addr_sel == 8'h75;
  assign mem_117_6_W0_addr = W0_addr[25:0];
  assign mem_117_6_W0_clk = W0_clk;
  assign mem_117_6_W0_data = W0_data[55:48];
  assign mem_117_6_W0_en = W0_en & W0_addr_sel == 8'h75;
  assign mem_117_6_W0_mask = W0_mask[6];
  assign mem_117_7_R0_addr = R0_addr[25:0];
  assign mem_117_7_R0_clk = R0_clk;
  assign mem_117_7_R0_en = R0_en & R0_addr_sel == 8'h75;
  assign mem_117_7_W0_addr = W0_addr[25:0];
  assign mem_117_7_W0_clk = W0_clk;
  assign mem_117_7_W0_data = W0_data[63:56];
  assign mem_117_7_W0_en = W0_en & W0_addr_sel == 8'h75;
  assign mem_117_7_W0_mask = W0_mask[7];
  assign mem_118_0_R0_addr = R0_addr[25:0];
  assign mem_118_0_R0_clk = R0_clk;
  assign mem_118_0_R0_en = R0_en & R0_addr_sel == 8'h76;
  assign mem_118_0_W0_addr = W0_addr[25:0];
  assign mem_118_0_W0_clk = W0_clk;
  assign mem_118_0_W0_data = W0_data[7:0];
  assign mem_118_0_W0_en = W0_en & W0_addr_sel == 8'h76;
  assign mem_118_0_W0_mask = W0_mask[0];
  assign mem_118_1_R0_addr = R0_addr[25:0];
  assign mem_118_1_R0_clk = R0_clk;
  assign mem_118_1_R0_en = R0_en & R0_addr_sel == 8'h76;
  assign mem_118_1_W0_addr = W0_addr[25:0];
  assign mem_118_1_W0_clk = W0_clk;
  assign mem_118_1_W0_data = W0_data[15:8];
  assign mem_118_1_W0_en = W0_en & W0_addr_sel == 8'h76;
  assign mem_118_1_W0_mask = W0_mask[1];
  assign mem_118_2_R0_addr = R0_addr[25:0];
  assign mem_118_2_R0_clk = R0_clk;
  assign mem_118_2_R0_en = R0_en & R0_addr_sel == 8'h76;
  assign mem_118_2_W0_addr = W0_addr[25:0];
  assign mem_118_2_W0_clk = W0_clk;
  assign mem_118_2_W0_data = W0_data[23:16];
  assign mem_118_2_W0_en = W0_en & W0_addr_sel == 8'h76;
  assign mem_118_2_W0_mask = W0_mask[2];
  assign mem_118_3_R0_addr = R0_addr[25:0];
  assign mem_118_3_R0_clk = R0_clk;
  assign mem_118_3_R0_en = R0_en & R0_addr_sel == 8'h76;
  assign mem_118_3_W0_addr = W0_addr[25:0];
  assign mem_118_3_W0_clk = W0_clk;
  assign mem_118_3_W0_data = W0_data[31:24];
  assign mem_118_3_W0_en = W0_en & W0_addr_sel == 8'h76;
  assign mem_118_3_W0_mask = W0_mask[3];
  assign mem_118_4_R0_addr = R0_addr[25:0];
  assign mem_118_4_R0_clk = R0_clk;
  assign mem_118_4_R0_en = R0_en & R0_addr_sel == 8'h76;
  assign mem_118_4_W0_addr = W0_addr[25:0];
  assign mem_118_4_W0_clk = W0_clk;
  assign mem_118_4_W0_data = W0_data[39:32];
  assign mem_118_4_W0_en = W0_en & W0_addr_sel == 8'h76;
  assign mem_118_4_W0_mask = W0_mask[4];
  assign mem_118_5_R0_addr = R0_addr[25:0];
  assign mem_118_5_R0_clk = R0_clk;
  assign mem_118_5_R0_en = R0_en & R0_addr_sel == 8'h76;
  assign mem_118_5_W0_addr = W0_addr[25:0];
  assign mem_118_5_W0_clk = W0_clk;
  assign mem_118_5_W0_data = W0_data[47:40];
  assign mem_118_5_W0_en = W0_en & W0_addr_sel == 8'h76;
  assign mem_118_5_W0_mask = W0_mask[5];
  assign mem_118_6_R0_addr = R0_addr[25:0];
  assign mem_118_6_R0_clk = R0_clk;
  assign mem_118_6_R0_en = R0_en & R0_addr_sel == 8'h76;
  assign mem_118_6_W0_addr = W0_addr[25:0];
  assign mem_118_6_W0_clk = W0_clk;
  assign mem_118_6_W0_data = W0_data[55:48];
  assign mem_118_6_W0_en = W0_en & W0_addr_sel == 8'h76;
  assign mem_118_6_W0_mask = W0_mask[6];
  assign mem_118_7_R0_addr = R0_addr[25:0];
  assign mem_118_7_R0_clk = R0_clk;
  assign mem_118_7_R0_en = R0_en & R0_addr_sel == 8'h76;
  assign mem_118_7_W0_addr = W0_addr[25:0];
  assign mem_118_7_W0_clk = W0_clk;
  assign mem_118_7_W0_data = W0_data[63:56];
  assign mem_118_7_W0_en = W0_en & W0_addr_sel == 8'h76;
  assign mem_118_7_W0_mask = W0_mask[7];
  assign mem_119_0_R0_addr = R0_addr[25:0];
  assign mem_119_0_R0_clk = R0_clk;
  assign mem_119_0_R0_en = R0_en & R0_addr_sel == 8'h77;
  assign mem_119_0_W0_addr = W0_addr[25:0];
  assign mem_119_0_W0_clk = W0_clk;
  assign mem_119_0_W0_data = W0_data[7:0];
  assign mem_119_0_W0_en = W0_en & W0_addr_sel == 8'h77;
  assign mem_119_0_W0_mask = W0_mask[0];
  assign mem_119_1_R0_addr = R0_addr[25:0];
  assign mem_119_1_R0_clk = R0_clk;
  assign mem_119_1_R0_en = R0_en & R0_addr_sel == 8'h77;
  assign mem_119_1_W0_addr = W0_addr[25:0];
  assign mem_119_1_W0_clk = W0_clk;
  assign mem_119_1_W0_data = W0_data[15:8];
  assign mem_119_1_W0_en = W0_en & W0_addr_sel == 8'h77;
  assign mem_119_1_W0_mask = W0_mask[1];
  assign mem_119_2_R0_addr = R0_addr[25:0];
  assign mem_119_2_R0_clk = R0_clk;
  assign mem_119_2_R0_en = R0_en & R0_addr_sel == 8'h77;
  assign mem_119_2_W0_addr = W0_addr[25:0];
  assign mem_119_2_W0_clk = W0_clk;
  assign mem_119_2_W0_data = W0_data[23:16];
  assign mem_119_2_W0_en = W0_en & W0_addr_sel == 8'h77;
  assign mem_119_2_W0_mask = W0_mask[2];
  assign mem_119_3_R0_addr = R0_addr[25:0];
  assign mem_119_3_R0_clk = R0_clk;
  assign mem_119_3_R0_en = R0_en & R0_addr_sel == 8'h77;
  assign mem_119_3_W0_addr = W0_addr[25:0];
  assign mem_119_3_W0_clk = W0_clk;
  assign mem_119_3_W0_data = W0_data[31:24];
  assign mem_119_3_W0_en = W0_en & W0_addr_sel == 8'h77;
  assign mem_119_3_W0_mask = W0_mask[3];
  assign mem_119_4_R0_addr = R0_addr[25:0];
  assign mem_119_4_R0_clk = R0_clk;
  assign mem_119_4_R0_en = R0_en & R0_addr_sel == 8'h77;
  assign mem_119_4_W0_addr = W0_addr[25:0];
  assign mem_119_4_W0_clk = W0_clk;
  assign mem_119_4_W0_data = W0_data[39:32];
  assign mem_119_4_W0_en = W0_en & W0_addr_sel == 8'h77;
  assign mem_119_4_W0_mask = W0_mask[4];
  assign mem_119_5_R0_addr = R0_addr[25:0];
  assign mem_119_5_R0_clk = R0_clk;
  assign mem_119_5_R0_en = R0_en & R0_addr_sel == 8'h77;
  assign mem_119_5_W0_addr = W0_addr[25:0];
  assign mem_119_5_W0_clk = W0_clk;
  assign mem_119_5_W0_data = W0_data[47:40];
  assign mem_119_5_W0_en = W0_en & W0_addr_sel == 8'h77;
  assign mem_119_5_W0_mask = W0_mask[5];
  assign mem_119_6_R0_addr = R0_addr[25:0];
  assign mem_119_6_R0_clk = R0_clk;
  assign mem_119_6_R0_en = R0_en & R0_addr_sel == 8'h77;
  assign mem_119_6_W0_addr = W0_addr[25:0];
  assign mem_119_6_W0_clk = W0_clk;
  assign mem_119_6_W0_data = W0_data[55:48];
  assign mem_119_6_W0_en = W0_en & W0_addr_sel == 8'h77;
  assign mem_119_6_W0_mask = W0_mask[6];
  assign mem_119_7_R0_addr = R0_addr[25:0];
  assign mem_119_7_R0_clk = R0_clk;
  assign mem_119_7_R0_en = R0_en & R0_addr_sel == 8'h77;
  assign mem_119_7_W0_addr = W0_addr[25:0];
  assign mem_119_7_W0_clk = W0_clk;
  assign mem_119_7_W0_data = W0_data[63:56];
  assign mem_119_7_W0_en = W0_en & W0_addr_sel == 8'h77;
  assign mem_119_7_W0_mask = W0_mask[7];
  assign mem_120_0_R0_addr = R0_addr[25:0];
  assign mem_120_0_R0_clk = R0_clk;
  assign mem_120_0_R0_en = R0_en & R0_addr_sel == 8'h78;
  assign mem_120_0_W0_addr = W0_addr[25:0];
  assign mem_120_0_W0_clk = W0_clk;
  assign mem_120_0_W0_data = W0_data[7:0];
  assign mem_120_0_W0_en = W0_en & W0_addr_sel == 8'h78;
  assign mem_120_0_W0_mask = W0_mask[0];
  assign mem_120_1_R0_addr = R0_addr[25:0];
  assign mem_120_1_R0_clk = R0_clk;
  assign mem_120_1_R0_en = R0_en & R0_addr_sel == 8'h78;
  assign mem_120_1_W0_addr = W0_addr[25:0];
  assign mem_120_1_W0_clk = W0_clk;
  assign mem_120_1_W0_data = W0_data[15:8];
  assign mem_120_1_W0_en = W0_en & W0_addr_sel == 8'h78;
  assign mem_120_1_W0_mask = W0_mask[1];
  assign mem_120_2_R0_addr = R0_addr[25:0];
  assign mem_120_2_R0_clk = R0_clk;
  assign mem_120_2_R0_en = R0_en & R0_addr_sel == 8'h78;
  assign mem_120_2_W0_addr = W0_addr[25:0];
  assign mem_120_2_W0_clk = W0_clk;
  assign mem_120_2_W0_data = W0_data[23:16];
  assign mem_120_2_W0_en = W0_en & W0_addr_sel == 8'h78;
  assign mem_120_2_W0_mask = W0_mask[2];
  assign mem_120_3_R0_addr = R0_addr[25:0];
  assign mem_120_3_R0_clk = R0_clk;
  assign mem_120_3_R0_en = R0_en & R0_addr_sel == 8'h78;
  assign mem_120_3_W0_addr = W0_addr[25:0];
  assign mem_120_3_W0_clk = W0_clk;
  assign mem_120_3_W0_data = W0_data[31:24];
  assign mem_120_3_W0_en = W0_en & W0_addr_sel == 8'h78;
  assign mem_120_3_W0_mask = W0_mask[3];
  assign mem_120_4_R0_addr = R0_addr[25:0];
  assign mem_120_4_R0_clk = R0_clk;
  assign mem_120_4_R0_en = R0_en & R0_addr_sel == 8'h78;
  assign mem_120_4_W0_addr = W0_addr[25:0];
  assign mem_120_4_W0_clk = W0_clk;
  assign mem_120_4_W0_data = W0_data[39:32];
  assign mem_120_4_W0_en = W0_en & W0_addr_sel == 8'h78;
  assign mem_120_4_W0_mask = W0_mask[4];
  assign mem_120_5_R0_addr = R0_addr[25:0];
  assign mem_120_5_R0_clk = R0_clk;
  assign mem_120_5_R0_en = R0_en & R0_addr_sel == 8'h78;
  assign mem_120_5_W0_addr = W0_addr[25:0];
  assign mem_120_5_W0_clk = W0_clk;
  assign mem_120_5_W0_data = W0_data[47:40];
  assign mem_120_5_W0_en = W0_en & W0_addr_sel == 8'h78;
  assign mem_120_5_W0_mask = W0_mask[5];
  assign mem_120_6_R0_addr = R0_addr[25:0];
  assign mem_120_6_R0_clk = R0_clk;
  assign mem_120_6_R0_en = R0_en & R0_addr_sel == 8'h78;
  assign mem_120_6_W0_addr = W0_addr[25:0];
  assign mem_120_6_W0_clk = W0_clk;
  assign mem_120_6_W0_data = W0_data[55:48];
  assign mem_120_6_W0_en = W0_en & W0_addr_sel == 8'h78;
  assign mem_120_6_W0_mask = W0_mask[6];
  assign mem_120_7_R0_addr = R0_addr[25:0];
  assign mem_120_7_R0_clk = R0_clk;
  assign mem_120_7_R0_en = R0_en & R0_addr_sel == 8'h78;
  assign mem_120_7_W0_addr = W0_addr[25:0];
  assign mem_120_7_W0_clk = W0_clk;
  assign mem_120_7_W0_data = W0_data[63:56];
  assign mem_120_7_W0_en = W0_en & W0_addr_sel == 8'h78;
  assign mem_120_7_W0_mask = W0_mask[7];
  assign mem_121_0_R0_addr = R0_addr[25:0];
  assign mem_121_0_R0_clk = R0_clk;
  assign mem_121_0_R0_en = R0_en & R0_addr_sel == 8'h79;
  assign mem_121_0_W0_addr = W0_addr[25:0];
  assign mem_121_0_W0_clk = W0_clk;
  assign mem_121_0_W0_data = W0_data[7:0];
  assign mem_121_0_W0_en = W0_en & W0_addr_sel == 8'h79;
  assign mem_121_0_W0_mask = W0_mask[0];
  assign mem_121_1_R0_addr = R0_addr[25:0];
  assign mem_121_1_R0_clk = R0_clk;
  assign mem_121_1_R0_en = R0_en & R0_addr_sel == 8'h79;
  assign mem_121_1_W0_addr = W0_addr[25:0];
  assign mem_121_1_W0_clk = W0_clk;
  assign mem_121_1_W0_data = W0_data[15:8];
  assign mem_121_1_W0_en = W0_en & W0_addr_sel == 8'h79;
  assign mem_121_1_W0_mask = W0_mask[1];
  assign mem_121_2_R0_addr = R0_addr[25:0];
  assign mem_121_2_R0_clk = R0_clk;
  assign mem_121_2_R0_en = R0_en & R0_addr_sel == 8'h79;
  assign mem_121_2_W0_addr = W0_addr[25:0];
  assign mem_121_2_W0_clk = W0_clk;
  assign mem_121_2_W0_data = W0_data[23:16];
  assign mem_121_2_W0_en = W0_en & W0_addr_sel == 8'h79;
  assign mem_121_2_W0_mask = W0_mask[2];
  assign mem_121_3_R0_addr = R0_addr[25:0];
  assign mem_121_3_R0_clk = R0_clk;
  assign mem_121_3_R0_en = R0_en & R0_addr_sel == 8'h79;
  assign mem_121_3_W0_addr = W0_addr[25:0];
  assign mem_121_3_W0_clk = W0_clk;
  assign mem_121_3_W0_data = W0_data[31:24];
  assign mem_121_3_W0_en = W0_en & W0_addr_sel == 8'h79;
  assign mem_121_3_W0_mask = W0_mask[3];
  assign mem_121_4_R0_addr = R0_addr[25:0];
  assign mem_121_4_R0_clk = R0_clk;
  assign mem_121_4_R0_en = R0_en & R0_addr_sel == 8'h79;
  assign mem_121_4_W0_addr = W0_addr[25:0];
  assign mem_121_4_W0_clk = W0_clk;
  assign mem_121_4_W0_data = W0_data[39:32];
  assign mem_121_4_W0_en = W0_en & W0_addr_sel == 8'h79;
  assign mem_121_4_W0_mask = W0_mask[4];
  assign mem_121_5_R0_addr = R0_addr[25:0];
  assign mem_121_5_R0_clk = R0_clk;
  assign mem_121_5_R0_en = R0_en & R0_addr_sel == 8'h79;
  assign mem_121_5_W0_addr = W0_addr[25:0];
  assign mem_121_5_W0_clk = W0_clk;
  assign mem_121_5_W0_data = W0_data[47:40];
  assign mem_121_5_W0_en = W0_en & W0_addr_sel == 8'h79;
  assign mem_121_5_W0_mask = W0_mask[5];
  assign mem_121_6_R0_addr = R0_addr[25:0];
  assign mem_121_6_R0_clk = R0_clk;
  assign mem_121_6_R0_en = R0_en & R0_addr_sel == 8'h79;
  assign mem_121_6_W0_addr = W0_addr[25:0];
  assign mem_121_6_W0_clk = W0_clk;
  assign mem_121_6_W0_data = W0_data[55:48];
  assign mem_121_6_W0_en = W0_en & W0_addr_sel == 8'h79;
  assign mem_121_6_W0_mask = W0_mask[6];
  assign mem_121_7_R0_addr = R0_addr[25:0];
  assign mem_121_7_R0_clk = R0_clk;
  assign mem_121_7_R0_en = R0_en & R0_addr_sel == 8'h79;
  assign mem_121_7_W0_addr = W0_addr[25:0];
  assign mem_121_7_W0_clk = W0_clk;
  assign mem_121_7_W0_data = W0_data[63:56];
  assign mem_121_7_W0_en = W0_en & W0_addr_sel == 8'h79;
  assign mem_121_7_W0_mask = W0_mask[7];
  assign mem_122_0_R0_addr = R0_addr[25:0];
  assign mem_122_0_R0_clk = R0_clk;
  assign mem_122_0_R0_en = R0_en & R0_addr_sel == 8'h7a;
  assign mem_122_0_W0_addr = W0_addr[25:0];
  assign mem_122_0_W0_clk = W0_clk;
  assign mem_122_0_W0_data = W0_data[7:0];
  assign mem_122_0_W0_en = W0_en & W0_addr_sel == 8'h7a;
  assign mem_122_0_W0_mask = W0_mask[0];
  assign mem_122_1_R0_addr = R0_addr[25:0];
  assign mem_122_1_R0_clk = R0_clk;
  assign mem_122_1_R0_en = R0_en & R0_addr_sel == 8'h7a;
  assign mem_122_1_W0_addr = W0_addr[25:0];
  assign mem_122_1_W0_clk = W0_clk;
  assign mem_122_1_W0_data = W0_data[15:8];
  assign mem_122_1_W0_en = W0_en & W0_addr_sel == 8'h7a;
  assign mem_122_1_W0_mask = W0_mask[1];
  assign mem_122_2_R0_addr = R0_addr[25:0];
  assign mem_122_2_R0_clk = R0_clk;
  assign mem_122_2_R0_en = R0_en & R0_addr_sel == 8'h7a;
  assign mem_122_2_W0_addr = W0_addr[25:0];
  assign mem_122_2_W0_clk = W0_clk;
  assign mem_122_2_W0_data = W0_data[23:16];
  assign mem_122_2_W0_en = W0_en & W0_addr_sel == 8'h7a;
  assign mem_122_2_W0_mask = W0_mask[2];
  assign mem_122_3_R0_addr = R0_addr[25:0];
  assign mem_122_3_R0_clk = R0_clk;
  assign mem_122_3_R0_en = R0_en & R0_addr_sel == 8'h7a;
  assign mem_122_3_W0_addr = W0_addr[25:0];
  assign mem_122_3_W0_clk = W0_clk;
  assign mem_122_3_W0_data = W0_data[31:24];
  assign mem_122_3_W0_en = W0_en & W0_addr_sel == 8'h7a;
  assign mem_122_3_W0_mask = W0_mask[3];
  assign mem_122_4_R0_addr = R0_addr[25:0];
  assign mem_122_4_R0_clk = R0_clk;
  assign mem_122_4_R0_en = R0_en & R0_addr_sel == 8'h7a;
  assign mem_122_4_W0_addr = W0_addr[25:0];
  assign mem_122_4_W0_clk = W0_clk;
  assign mem_122_4_W0_data = W0_data[39:32];
  assign mem_122_4_W0_en = W0_en & W0_addr_sel == 8'h7a;
  assign mem_122_4_W0_mask = W0_mask[4];
  assign mem_122_5_R0_addr = R0_addr[25:0];
  assign mem_122_5_R0_clk = R0_clk;
  assign mem_122_5_R0_en = R0_en & R0_addr_sel == 8'h7a;
  assign mem_122_5_W0_addr = W0_addr[25:0];
  assign mem_122_5_W0_clk = W0_clk;
  assign mem_122_5_W0_data = W0_data[47:40];
  assign mem_122_5_W0_en = W0_en & W0_addr_sel == 8'h7a;
  assign mem_122_5_W0_mask = W0_mask[5];
  assign mem_122_6_R0_addr = R0_addr[25:0];
  assign mem_122_6_R0_clk = R0_clk;
  assign mem_122_6_R0_en = R0_en & R0_addr_sel == 8'h7a;
  assign mem_122_6_W0_addr = W0_addr[25:0];
  assign mem_122_6_W0_clk = W0_clk;
  assign mem_122_6_W0_data = W0_data[55:48];
  assign mem_122_6_W0_en = W0_en & W0_addr_sel == 8'h7a;
  assign mem_122_6_W0_mask = W0_mask[6];
  assign mem_122_7_R0_addr = R0_addr[25:0];
  assign mem_122_7_R0_clk = R0_clk;
  assign mem_122_7_R0_en = R0_en & R0_addr_sel == 8'h7a;
  assign mem_122_7_W0_addr = W0_addr[25:0];
  assign mem_122_7_W0_clk = W0_clk;
  assign mem_122_7_W0_data = W0_data[63:56];
  assign mem_122_7_W0_en = W0_en & W0_addr_sel == 8'h7a;
  assign mem_122_7_W0_mask = W0_mask[7];
  assign mem_123_0_R0_addr = R0_addr[25:0];
  assign mem_123_0_R0_clk = R0_clk;
  assign mem_123_0_R0_en = R0_en & R0_addr_sel == 8'h7b;
  assign mem_123_0_W0_addr = W0_addr[25:0];
  assign mem_123_0_W0_clk = W0_clk;
  assign mem_123_0_W0_data = W0_data[7:0];
  assign mem_123_0_W0_en = W0_en & W0_addr_sel == 8'h7b;
  assign mem_123_0_W0_mask = W0_mask[0];
  assign mem_123_1_R0_addr = R0_addr[25:0];
  assign mem_123_1_R0_clk = R0_clk;
  assign mem_123_1_R0_en = R0_en & R0_addr_sel == 8'h7b;
  assign mem_123_1_W0_addr = W0_addr[25:0];
  assign mem_123_1_W0_clk = W0_clk;
  assign mem_123_1_W0_data = W0_data[15:8];
  assign mem_123_1_W0_en = W0_en & W0_addr_sel == 8'h7b;
  assign mem_123_1_W0_mask = W0_mask[1];
  assign mem_123_2_R0_addr = R0_addr[25:0];
  assign mem_123_2_R0_clk = R0_clk;
  assign mem_123_2_R0_en = R0_en & R0_addr_sel == 8'h7b;
  assign mem_123_2_W0_addr = W0_addr[25:0];
  assign mem_123_2_W0_clk = W0_clk;
  assign mem_123_2_W0_data = W0_data[23:16];
  assign mem_123_2_W0_en = W0_en & W0_addr_sel == 8'h7b;
  assign mem_123_2_W0_mask = W0_mask[2];
  assign mem_123_3_R0_addr = R0_addr[25:0];
  assign mem_123_3_R0_clk = R0_clk;
  assign mem_123_3_R0_en = R0_en & R0_addr_sel == 8'h7b;
  assign mem_123_3_W0_addr = W0_addr[25:0];
  assign mem_123_3_W0_clk = W0_clk;
  assign mem_123_3_W0_data = W0_data[31:24];
  assign mem_123_3_W0_en = W0_en & W0_addr_sel == 8'h7b;
  assign mem_123_3_W0_mask = W0_mask[3];
  assign mem_123_4_R0_addr = R0_addr[25:0];
  assign mem_123_4_R0_clk = R0_clk;
  assign mem_123_4_R0_en = R0_en & R0_addr_sel == 8'h7b;
  assign mem_123_4_W0_addr = W0_addr[25:0];
  assign mem_123_4_W0_clk = W0_clk;
  assign mem_123_4_W0_data = W0_data[39:32];
  assign mem_123_4_W0_en = W0_en & W0_addr_sel == 8'h7b;
  assign mem_123_4_W0_mask = W0_mask[4];
  assign mem_123_5_R0_addr = R0_addr[25:0];
  assign mem_123_5_R0_clk = R0_clk;
  assign mem_123_5_R0_en = R0_en & R0_addr_sel == 8'h7b;
  assign mem_123_5_W0_addr = W0_addr[25:0];
  assign mem_123_5_W0_clk = W0_clk;
  assign mem_123_5_W0_data = W0_data[47:40];
  assign mem_123_5_W0_en = W0_en & W0_addr_sel == 8'h7b;
  assign mem_123_5_W0_mask = W0_mask[5];
  assign mem_123_6_R0_addr = R0_addr[25:0];
  assign mem_123_6_R0_clk = R0_clk;
  assign mem_123_6_R0_en = R0_en & R0_addr_sel == 8'h7b;
  assign mem_123_6_W0_addr = W0_addr[25:0];
  assign mem_123_6_W0_clk = W0_clk;
  assign mem_123_6_W0_data = W0_data[55:48];
  assign mem_123_6_W0_en = W0_en & W0_addr_sel == 8'h7b;
  assign mem_123_6_W0_mask = W0_mask[6];
  assign mem_123_7_R0_addr = R0_addr[25:0];
  assign mem_123_7_R0_clk = R0_clk;
  assign mem_123_7_R0_en = R0_en & R0_addr_sel == 8'h7b;
  assign mem_123_7_W0_addr = W0_addr[25:0];
  assign mem_123_7_W0_clk = W0_clk;
  assign mem_123_7_W0_data = W0_data[63:56];
  assign mem_123_7_W0_en = W0_en & W0_addr_sel == 8'h7b;
  assign mem_123_7_W0_mask = W0_mask[7];
  assign mem_124_0_R0_addr = R0_addr[25:0];
  assign mem_124_0_R0_clk = R0_clk;
  assign mem_124_0_R0_en = R0_en & R0_addr_sel == 8'h7c;
  assign mem_124_0_W0_addr = W0_addr[25:0];
  assign mem_124_0_W0_clk = W0_clk;
  assign mem_124_0_W0_data = W0_data[7:0];
  assign mem_124_0_W0_en = W0_en & W0_addr_sel == 8'h7c;
  assign mem_124_0_W0_mask = W0_mask[0];
  assign mem_124_1_R0_addr = R0_addr[25:0];
  assign mem_124_1_R0_clk = R0_clk;
  assign mem_124_1_R0_en = R0_en & R0_addr_sel == 8'h7c;
  assign mem_124_1_W0_addr = W0_addr[25:0];
  assign mem_124_1_W0_clk = W0_clk;
  assign mem_124_1_W0_data = W0_data[15:8];
  assign mem_124_1_W0_en = W0_en & W0_addr_sel == 8'h7c;
  assign mem_124_1_W0_mask = W0_mask[1];
  assign mem_124_2_R0_addr = R0_addr[25:0];
  assign mem_124_2_R0_clk = R0_clk;
  assign mem_124_2_R0_en = R0_en & R0_addr_sel == 8'h7c;
  assign mem_124_2_W0_addr = W0_addr[25:0];
  assign mem_124_2_W0_clk = W0_clk;
  assign mem_124_2_W0_data = W0_data[23:16];
  assign mem_124_2_W0_en = W0_en & W0_addr_sel == 8'h7c;
  assign mem_124_2_W0_mask = W0_mask[2];
  assign mem_124_3_R0_addr = R0_addr[25:0];
  assign mem_124_3_R0_clk = R0_clk;
  assign mem_124_3_R0_en = R0_en & R0_addr_sel == 8'h7c;
  assign mem_124_3_W0_addr = W0_addr[25:0];
  assign mem_124_3_W0_clk = W0_clk;
  assign mem_124_3_W0_data = W0_data[31:24];
  assign mem_124_3_W0_en = W0_en & W0_addr_sel == 8'h7c;
  assign mem_124_3_W0_mask = W0_mask[3];
  assign mem_124_4_R0_addr = R0_addr[25:0];
  assign mem_124_4_R0_clk = R0_clk;
  assign mem_124_4_R0_en = R0_en & R0_addr_sel == 8'h7c;
  assign mem_124_4_W0_addr = W0_addr[25:0];
  assign mem_124_4_W0_clk = W0_clk;
  assign mem_124_4_W0_data = W0_data[39:32];
  assign mem_124_4_W0_en = W0_en & W0_addr_sel == 8'h7c;
  assign mem_124_4_W0_mask = W0_mask[4];
  assign mem_124_5_R0_addr = R0_addr[25:0];
  assign mem_124_5_R0_clk = R0_clk;
  assign mem_124_5_R0_en = R0_en & R0_addr_sel == 8'h7c;
  assign mem_124_5_W0_addr = W0_addr[25:0];
  assign mem_124_5_W0_clk = W0_clk;
  assign mem_124_5_W0_data = W0_data[47:40];
  assign mem_124_5_W0_en = W0_en & W0_addr_sel == 8'h7c;
  assign mem_124_5_W0_mask = W0_mask[5];
  assign mem_124_6_R0_addr = R0_addr[25:0];
  assign mem_124_6_R0_clk = R0_clk;
  assign mem_124_6_R0_en = R0_en & R0_addr_sel == 8'h7c;
  assign mem_124_6_W0_addr = W0_addr[25:0];
  assign mem_124_6_W0_clk = W0_clk;
  assign mem_124_6_W0_data = W0_data[55:48];
  assign mem_124_6_W0_en = W0_en & W0_addr_sel == 8'h7c;
  assign mem_124_6_W0_mask = W0_mask[6];
  assign mem_124_7_R0_addr = R0_addr[25:0];
  assign mem_124_7_R0_clk = R0_clk;
  assign mem_124_7_R0_en = R0_en & R0_addr_sel == 8'h7c;
  assign mem_124_7_W0_addr = W0_addr[25:0];
  assign mem_124_7_W0_clk = W0_clk;
  assign mem_124_7_W0_data = W0_data[63:56];
  assign mem_124_7_W0_en = W0_en & W0_addr_sel == 8'h7c;
  assign mem_124_7_W0_mask = W0_mask[7];
  assign mem_125_0_R0_addr = R0_addr[25:0];
  assign mem_125_0_R0_clk = R0_clk;
  assign mem_125_0_R0_en = R0_en & R0_addr_sel == 8'h7d;
  assign mem_125_0_W0_addr = W0_addr[25:0];
  assign mem_125_0_W0_clk = W0_clk;
  assign mem_125_0_W0_data = W0_data[7:0];
  assign mem_125_0_W0_en = W0_en & W0_addr_sel == 8'h7d;
  assign mem_125_0_W0_mask = W0_mask[0];
  assign mem_125_1_R0_addr = R0_addr[25:0];
  assign mem_125_1_R0_clk = R0_clk;
  assign mem_125_1_R0_en = R0_en & R0_addr_sel == 8'h7d;
  assign mem_125_1_W0_addr = W0_addr[25:0];
  assign mem_125_1_W0_clk = W0_clk;
  assign mem_125_1_W0_data = W0_data[15:8];
  assign mem_125_1_W0_en = W0_en & W0_addr_sel == 8'h7d;
  assign mem_125_1_W0_mask = W0_mask[1];
  assign mem_125_2_R0_addr = R0_addr[25:0];
  assign mem_125_2_R0_clk = R0_clk;
  assign mem_125_2_R0_en = R0_en & R0_addr_sel == 8'h7d;
  assign mem_125_2_W0_addr = W0_addr[25:0];
  assign mem_125_2_W0_clk = W0_clk;
  assign mem_125_2_W0_data = W0_data[23:16];
  assign mem_125_2_W0_en = W0_en & W0_addr_sel == 8'h7d;
  assign mem_125_2_W0_mask = W0_mask[2];
  assign mem_125_3_R0_addr = R0_addr[25:0];
  assign mem_125_3_R0_clk = R0_clk;
  assign mem_125_3_R0_en = R0_en & R0_addr_sel == 8'h7d;
  assign mem_125_3_W0_addr = W0_addr[25:0];
  assign mem_125_3_W0_clk = W0_clk;
  assign mem_125_3_W0_data = W0_data[31:24];
  assign mem_125_3_W0_en = W0_en & W0_addr_sel == 8'h7d;
  assign mem_125_3_W0_mask = W0_mask[3];
  assign mem_125_4_R0_addr = R0_addr[25:0];
  assign mem_125_4_R0_clk = R0_clk;
  assign mem_125_4_R0_en = R0_en & R0_addr_sel == 8'h7d;
  assign mem_125_4_W0_addr = W0_addr[25:0];
  assign mem_125_4_W0_clk = W0_clk;
  assign mem_125_4_W0_data = W0_data[39:32];
  assign mem_125_4_W0_en = W0_en & W0_addr_sel == 8'h7d;
  assign mem_125_4_W0_mask = W0_mask[4];
  assign mem_125_5_R0_addr = R0_addr[25:0];
  assign mem_125_5_R0_clk = R0_clk;
  assign mem_125_5_R0_en = R0_en & R0_addr_sel == 8'h7d;
  assign mem_125_5_W0_addr = W0_addr[25:0];
  assign mem_125_5_W0_clk = W0_clk;
  assign mem_125_5_W0_data = W0_data[47:40];
  assign mem_125_5_W0_en = W0_en & W0_addr_sel == 8'h7d;
  assign mem_125_5_W0_mask = W0_mask[5];
  assign mem_125_6_R0_addr = R0_addr[25:0];
  assign mem_125_6_R0_clk = R0_clk;
  assign mem_125_6_R0_en = R0_en & R0_addr_sel == 8'h7d;
  assign mem_125_6_W0_addr = W0_addr[25:0];
  assign mem_125_6_W0_clk = W0_clk;
  assign mem_125_6_W0_data = W0_data[55:48];
  assign mem_125_6_W0_en = W0_en & W0_addr_sel == 8'h7d;
  assign mem_125_6_W0_mask = W0_mask[6];
  assign mem_125_7_R0_addr = R0_addr[25:0];
  assign mem_125_7_R0_clk = R0_clk;
  assign mem_125_7_R0_en = R0_en & R0_addr_sel == 8'h7d;
  assign mem_125_7_W0_addr = W0_addr[25:0];
  assign mem_125_7_W0_clk = W0_clk;
  assign mem_125_7_W0_data = W0_data[63:56];
  assign mem_125_7_W0_en = W0_en & W0_addr_sel == 8'h7d;
  assign mem_125_7_W0_mask = W0_mask[7];
  assign mem_126_0_R0_addr = R0_addr[25:0];
  assign mem_126_0_R0_clk = R0_clk;
  assign mem_126_0_R0_en = R0_en & R0_addr_sel == 8'h7e;
  assign mem_126_0_W0_addr = W0_addr[25:0];
  assign mem_126_0_W0_clk = W0_clk;
  assign mem_126_0_W0_data = W0_data[7:0];
  assign mem_126_0_W0_en = W0_en & W0_addr_sel == 8'h7e;
  assign mem_126_0_W0_mask = W0_mask[0];
  assign mem_126_1_R0_addr = R0_addr[25:0];
  assign mem_126_1_R0_clk = R0_clk;
  assign mem_126_1_R0_en = R0_en & R0_addr_sel == 8'h7e;
  assign mem_126_1_W0_addr = W0_addr[25:0];
  assign mem_126_1_W0_clk = W0_clk;
  assign mem_126_1_W0_data = W0_data[15:8];
  assign mem_126_1_W0_en = W0_en & W0_addr_sel == 8'h7e;
  assign mem_126_1_W0_mask = W0_mask[1];
  assign mem_126_2_R0_addr = R0_addr[25:0];
  assign mem_126_2_R0_clk = R0_clk;
  assign mem_126_2_R0_en = R0_en & R0_addr_sel == 8'h7e;
  assign mem_126_2_W0_addr = W0_addr[25:0];
  assign mem_126_2_W0_clk = W0_clk;
  assign mem_126_2_W0_data = W0_data[23:16];
  assign mem_126_2_W0_en = W0_en & W0_addr_sel == 8'h7e;
  assign mem_126_2_W0_mask = W0_mask[2];
  assign mem_126_3_R0_addr = R0_addr[25:0];
  assign mem_126_3_R0_clk = R0_clk;
  assign mem_126_3_R0_en = R0_en & R0_addr_sel == 8'h7e;
  assign mem_126_3_W0_addr = W0_addr[25:0];
  assign mem_126_3_W0_clk = W0_clk;
  assign mem_126_3_W0_data = W0_data[31:24];
  assign mem_126_3_W0_en = W0_en & W0_addr_sel == 8'h7e;
  assign mem_126_3_W0_mask = W0_mask[3];
  assign mem_126_4_R0_addr = R0_addr[25:0];
  assign mem_126_4_R0_clk = R0_clk;
  assign mem_126_4_R0_en = R0_en & R0_addr_sel == 8'h7e;
  assign mem_126_4_W0_addr = W0_addr[25:0];
  assign mem_126_4_W0_clk = W0_clk;
  assign mem_126_4_W0_data = W0_data[39:32];
  assign mem_126_4_W0_en = W0_en & W0_addr_sel == 8'h7e;
  assign mem_126_4_W0_mask = W0_mask[4];
  assign mem_126_5_R0_addr = R0_addr[25:0];
  assign mem_126_5_R0_clk = R0_clk;
  assign mem_126_5_R0_en = R0_en & R0_addr_sel == 8'h7e;
  assign mem_126_5_W0_addr = W0_addr[25:0];
  assign mem_126_5_W0_clk = W0_clk;
  assign mem_126_5_W0_data = W0_data[47:40];
  assign mem_126_5_W0_en = W0_en & W0_addr_sel == 8'h7e;
  assign mem_126_5_W0_mask = W0_mask[5];
  assign mem_126_6_R0_addr = R0_addr[25:0];
  assign mem_126_6_R0_clk = R0_clk;
  assign mem_126_6_R0_en = R0_en & R0_addr_sel == 8'h7e;
  assign mem_126_6_W0_addr = W0_addr[25:0];
  assign mem_126_6_W0_clk = W0_clk;
  assign mem_126_6_W0_data = W0_data[55:48];
  assign mem_126_6_W0_en = W0_en & W0_addr_sel == 8'h7e;
  assign mem_126_6_W0_mask = W0_mask[6];
  assign mem_126_7_R0_addr = R0_addr[25:0];
  assign mem_126_7_R0_clk = R0_clk;
  assign mem_126_7_R0_en = R0_en & R0_addr_sel == 8'h7e;
  assign mem_126_7_W0_addr = W0_addr[25:0];
  assign mem_126_7_W0_clk = W0_clk;
  assign mem_126_7_W0_data = W0_data[63:56];
  assign mem_126_7_W0_en = W0_en & W0_addr_sel == 8'h7e;
  assign mem_126_7_W0_mask = W0_mask[7];
  assign mem_127_0_R0_addr = R0_addr[25:0];
  assign mem_127_0_R0_clk = R0_clk;
  assign mem_127_0_R0_en = R0_en & R0_addr_sel == 8'h7f;
  assign mem_127_0_W0_addr = W0_addr[25:0];
  assign mem_127_0_W0_clk = W0_clk;
  assign mem_127_0_W0_data = W0_data[7:0];
  assign mem_127_0_W0_en = W0_en & W0_addr_sel == 8'h7f;
  assign mem_127_0_W0_mask = W0_mask[0];
  assign mem_127_1_R0_addr = R0_addr[25:0];
  assign mem_127_1_R0_clk = R0_clk;
  assign mem_127_1_R0_en = R0_en & R0_addr_sel == 8'h7f;
  assign mem_127_1_W0_addr = W0_addr[25:0];
  assign mem_127_1_W0_clk = W0_clk;
  assign mem_127_1_W0_data = W0_data[15:8];
  assign mem_127_1_W0_en = W0_en & W0_addr_sel == 8'h7f;
  assign mem_127_1_W0_mask = W0_mask[1];
  assign mem_127_2_R0_addr = R0_addr[25:0];
  assign mem_127_2_R0_clk = R0_clk;
  assign mem_127_2_R0_en = R0_en & R0_addr_sel == 8'h7f;
  assign mem_127_2_W0_addr = W0_addr[25:0];
  assign mem_127_2_W0_clk = W0_clk;
  assign mem_127_2_W0_data = W0_data[23:16];
  assign mem_127_2_W0_en = W0_en & W0_addr_sel == 8'h7f;
  assign mem_127_2_W0_mask = W0_mask[2];
  assign mem_127_3_R0_addr = R0_addr[25:0];
  assign mem_127_3_R0_clk = R0_clk;
  assign mem_127_3_R0_en = R0_en & R0_addr_sel == 8'h7f;
  assign mem_127_3_W0_addr = W0_addr[25:0];
  assign mem_127_3_W0_clk = W0_clk;
  assign mem_127_3_W0_data = W0_data[31:24];
  assign mem_127_3_W0_en = W0_en & W0_addr_sel == 8'h7f;
  assign mem_127_3_W0_mask = W0_mask[3];
  assign mem_127_4_R0_addr = R0_addr[25:0];
  assign mem_127_4_R0_clk = R0_clk;
  assign mem_127_4_R0_en = R0_en & R0_addr_sel == 8'h7f;
  assign mem_127_4_W0_addr = W0_addr[25:0];
  assign mem_127_4_W0_clk = W0_clk;
  assign mem_127_4_W0_data = W0_data[39:32];
  assign mem_127_4_W0_en = W0_en & W0_addr_sel == 8'h7f;
  assign mem_127_4_W0_mask = W0_mask[4];
  assign mem_127_5_R0_addr = R0_addr[25:0];
  assign mem_127_5_R0_clk = R0_clk;
  assign mem_127_5_R0_en = R0_en & R0_addr_sel == 8'h7f;
  assign mem_127_5_W0_addr = W0_addr[25:0];
  assign mem_127_5_W0_clk = W0_clk;
  assign mem_127_5_W0_data = W0_data[47:40];
  assign mem_127_5_W0_en = W0_en & W0_addr_sel == 8'h7f;
  assign mem_127_5_W0_mask = W0_mask[5];
  assign mem_127_6_R0_addr = R0_addr[25:0];
  assign mem_127_6_R0_clk = R0_clk;
  assign mem_127_6_R0_en = R0_en & R0_addr_sel == 8'h7f;
  assign mem_127_6_W0_addr = W0_addr[25:0];
  assign mem_127_6_W0_clk = W0_clk;
  assign mem_127_6_W0_data = W0_data[55:48];
  assign mem_127_6_W0_en = W0_en & W0_addr_sel == 8'h7f;
  assign mem_127_6_W0_mask = W0_mask[6];
  assign mem_127_7_R0_addr = R0_addr[25:0];
  assign mem_127_7_R0_clk = R0_clk;
  assign mem_127_7_R0_en = R0_en & R0_addr_sel == 8'h7f;
  assign mem_127_7_W0_addr = W0_addr[25:0];
  assign mem_127_7_W0_clk = W0_clk;
  assign mem_127_7_W0_data = W0_data[63:56];
  assign mem_127_7_W0_en = W0_en & W0_addr_sel == 8'h7f;
  assign mem_127_7_W0_mask = W0_mask[7];
  assign mem_128_0_R0_addr = R0_addr[25:0];
  assign mem_128_0_R0_clk = R0_clk;
  assign mem_128_0_R0_en = R0_en & R0_addr_sel == 8'h80;
  assign mem_128_0_W0_addr = W0_addr[25:0];
  assign mem_128_0_W0_clk = W0_clk;
  assign mem_128_0_W0_data = W0_data[7:0];
  assign mem_128_0_W0_en = W0_en & W0_addr_sel == 8'h80;
  assign mem_128_0_W0_mask = W0_mask[0];
  assign mem_128_1_R0_addr = R0_addr[25:0];
  assign mem_128_1_R0_clk = R0_clk;
  assign mem_128_1_R0_en = R0_en & R0_addr_sel == 8'h80;
  assign mem_128_1_W0_addr = W0_addr[25:0];
  assign mem_128_1_W0_clk = W0_clk;
  assign mem_128_1_W0_data = W0_data[15:8];
  assign mem_128_1_W0_en = W0_en & W0_addr_sel == 8'h80;
  assign mem_128_1_W0_mask = W0_mask[1];
  assign mem_128_2_R0_addr = R0_addr[25:0];
  assign mem_128_2_R0_clk = R0_clk;
  assign mem_128_2_R0_en = R0_en & R0_addr_sel == 8'h80;
  assign mem_128_2_W0_addr = W0_addr[25:0];
  assign mem_128_2_W0_clk = W0_clk;
  assign mem_128_2_W0_data = W0_data[23:16];
  assign mem_128_2_W0_en = W0_en & W0_addr_sel == 8'h80;
  assign mem_128_2_W0_mask = W0_mask[2];
  assign mem_128_3_R0_addr = R0_addr[25:0];
  assign mem_128_3_R0_clk = R0_clk;
  assign mem_128_3_R0_en = R0_en & R0_addr_sel == 8'h80;
  assign mem_128_3_W0_addr = W0_addr[25:0];
  assign mem_128_3_W0_clk = W0_clk;
  assign mem_128_3_W0_data = W0_data[31:24];
  assign mem_128_3_W0_en = W0_en & W0_addr_sel == 8'h80;
  assign mem_128_3_W0_mask = W0_mask[3];
  assign mem_128_4_R0_addr = R0_addr[25:0];
  assign mem_128_4_R0_clk = R0_clk;
  assign mem_128_4_R0_en = R0_en & R0_addr_sel == 8'h80;
  assign mem_128_4_W0_addr = W0_addr[25:0];
  assign mem_128_4_W0_clk = W0_clk;
  assign mem_128_4_W0_data = W0_data[39:32];
  assign mem_128_4_W0_en = W0_en & W0_addr_sel == 8'h80;
  assign mem_128_4_W0_mask = W0_mask[4];
  assign mem_128_5_R0_addr = R0_addr[25:0];
  assign mem_128_5_R0_clk = R0_clk;
  assign mem_128_5_R0_en = R0_en & R0_addr_sel == 8'h80;
  assign mem_128_5_W0_addr = W0_addr[25:0];
  assign mem_128_5_W0_clk = W0_clk;
  assign mem_128_5_W0_data = W0_data[47:40];
  assign mem_128_5_W0_en = W0_en & W0_addr_sel == 8'h80;
  assign mem_128_5_W0_mask = W0_mask[5];
  assign mem_128_6_R0_addr = R0_addr[25:0];
  assign mem_128_6_R0_clk = R0_clk;
  assign mem_128_6_R0_en = R0_en & R0_addr_sel == 8'h80;
  assign mem_128_6_W0_addr = W0_addr[25:0];
  assign mem_128_6_W0_clk = W0_clk;
  assign mem_128_6_W0_data = W0_data[55:48];
  assign mem_128_6_W0_en = W0_en & W0_addr_sel == 8'h80;
  assign mem_128_6_W0_mask = W0_mask[6];
  assign mem_128_7_R0_addr = R0_addr[25:0];
  assign mem_128_7_R0_clk = R0_clk;
  assign mem_128_7_R0_en = R0_en & R0_addr_sel == 8'h80;
  assign mem_128_7_W0_addr = W0_addr[25:0];
  assign mem_128_7_W0_clk = W0_clk;
  assign mem_128_7_W0_data = W0_data[63:56];
  assign mem_128_7_W0_en = W0_en & W0_addr_sel == 8'h80;
  assign mem_128_7_W0_mask = W0_mask[7];
  assign mem_129_0_R0_addr = R0_addr[25:0];
  assign mem_129_0_R0_clk = R0_clk;
  assign mem_129_0_R0_en = R0_en & R0_addr_sel == 8'h81;
  assign mem_129_0_W0_addr = W0_addr[25:0];
  assign mem_129_0_W0_clk = W0_clk;
  assign mem_129_0_W0_data = W0_data[7:0];
  assign mem_129_0_W0_en = W0_en & W0_addr_sel == 8'h81;
  assign mem_129_0_W0_mask = W0_mask[0];
  assign mem_129_1_R0_addr = R0_addr[25:0];
  assign mem_129_1_R0_clk = R0_clk;
  assign mem_129_1_R0_en = R0_en & R0_addr_sel == 8'h81;
  assign mem_129_1_W0_addr = W0_addr[25:0];
  assign mem_129_1_W0_clk = W0_clk;
  assign mem_129_1_W0_data = W0_data[15:8];
  assign mem_129_1_W0_en = W0_en & W0_addr_sel == 8'h81;
  assign mem_129_1_W0_mask = W0_mask[1];
  assign mem_129_2_R0_addr = R0_addr[25:0];
  assign mem_129_2_R0_clk = R0_clk;
  assign mem_129_2_R0_en = R0_en & R0_addr_sel == 8'h81;
  assign mem_129_2_W0_addr = W0_addr[25:0];
  assign mem_129_2_W0_clk = W0_clk;
  assign mem_129_2_W0_data = W0_data[23:16];
  assign mem_129_2_W0_en = W0_en & W0_addr_sel == 8'h81;
  assign mem_129_2_W0_mask = W0_mask[2];
  assign mem_129_3_R0_addr = R0_addr[25:0];
  assign mem_129_3_R0_clk = R0_clk;
  assign mem_129_3_R0_en = R0_en & R0_addr_sel == 8'h81;
  assign mem_129_3_W0_addr = W0_addr[25:0];
  assign mem_129_3_W0_clk = W0_clk;
  assign mem_129_3_W0_data = W0_data[31:24];
  assign mem_129_3_W0_en = W0_en & W0_addr_sel == 8'h81;
  assign mem_129_3_W0_mask = W0_mask[3];
  assign mem_129_4_R0_addr = R0_addr[25:0];
  assign mem_129_4_R0_clk = R0_clk;
  assign mem_129_4_R0_en = R0_en & R0_addr_sel == 8'h81;
  assign mem_129_4_W0_addr = W0_addr[25:0];
  assign mem_129_4_W0_clk = W0_clk;
  assign mem_129_4_W0_data = W0_data[39:32];
  assign mem_129_4_W0_en = W0_en & W0_addr_sel == 8'h81;
  assign mem_129_4_W0_mask = W0_mask[4];
  assign mem_129_5_R0_addr = R0_addr[25:0];
  assign mem_129_5_R0_clk = R0_clk;
  assign mem_129_5_R0_en = R0_en & R0_addr_sel == 8'h81;
  assign mem_129_5_W0_addr = W0_addr[25:0];
  assign mem_129_5_W0_clk = W0_clk;
  assign mem_129_5_W0_data = W0_data[47:40];
  assign mem_129_5_W0_en = W0_en & W0_addr_sel == 8'h81;
  assign mem_129_5_W0_mask = W0_mask[5];
  assign mem_129_6_R0_addr = R0_addr[25:0];
  assign mem_129_6_R0_clk = R0_clk;
  assign mem_129_6_R0_en = R0_en & R0_addr_sel == 8'h81;
  assign mem_129_6_W0_addr = W0_addr[25:0];
  assign mem_129_6_W0_clk = W0_clk;
  assign mem_129_6_W0_data = W0_data[55:48];
  assign mem_129_6_W0_en = W0_en & W0_addr_sel == 8'h81;
  assign mem_129_6_W0_mask = W0_mask[6];
  assign mem_129_7_R0_addr = R0_addr[25:0];
  assign mem_129_7_R0_clk = R0_clk;
  assign mem_129_7_R0_en = R0_en & R0_addr_sel == 8'h81;
  assign mem_129_7_W0_addr = W0_addr[25:0];
  assign mem_129_7_W0_clk = W0_clk;
  assign mem_129_7_W0_data = W0_data[63:56];
  assign mem_129_7_W0_en = W0_en & W0_addr_sel == 8'h81;
  assign mem_129_7_W0_mask = W0_mask[7];
  assign mem_130_0_R0_addr = R0_addr[25:0];
  assign mem_130_0_R0_clk = R0_clk;
  assign mem_130_0_R0_en = R0_en & R0_addr_sel == 8'h82;
  assign mem_130_0_W0_addr = W0_addr[25:0];
  assign mem_130_0_W0_clk = W0_clk;
  assign mem_130_0_W0_data = W0_data[7:0];
  assign mem_130_0_W0_en = W0_en & W0_addr_sel == 8'h82;
  assign mem_130_0_W0_mask = W0_mask[0];
  assign mem_130_1_R0_addr = R0_addr[25:0];
  assign mem_130_1_R0_clk = R0_clk;
  assign mem_130_1_R0_en = R0_en & R0_addr_sel == 8'h82;
  assign mem_130_1_W0_addr = W0_addr[25:0];
  assign mem_130_1_W0_clk = W0_clk;
  assign mem_130_1_W0_data = W0_data[15:8];
  assign mem_130_1_W0_en = W0_en & W0_addr_sel == 8'h82;
  assign mem_130_1_W0_mask = W0_mask[1];
  assign mem_130_2_R0_addr = R0_addr[25:0];
  assign mem_130_2_R0_clk = R0_clk;
  assign mem_130_2_R0_en = R0_en & R0_addr_sel == 8'h82;
  assign mem_130_2_W0_addr = W0_addr[25:0];
  assign mem_130_2_W0_clk = W0_clk;
  assign mem_130_2_W0_data = W0_data[23:16];
  assign mem_130_2_W0_en = W0_en & W0_addr_sel == 8'h82;
  assign mem_130_2_W0_mask = W0_mask[2];
  assign mem_130_3_R0_addr = R0_addr[25:0];
  assign mem_130_3_R0_clk = R0_clk;
  assign mem_130_3_R0_en = R0_en & R0_addr_sel == 8'h82;
  assign mem_130_3_W0_addr = W0_addr[25:0];
  assign mem_130_3_W0_clk = W0_clk;
  assign mem_130_3_W0_data = W0_data[31:24];
  assign mem_130_3_W0_en = W0_en & W0_addr_sel == 8'h82;
  assign mem_130_3_W0_mask = W0_mask[3];
  assign mem_130_4_R0_addr = R0_addr[25:0];
  assign mem_130_4_R0_clk = R0_clk;
  assign mem_130_4_R0_en = R0_en & R0_addr_sel == 8'h82;
  assign mem_130_4_W0_addr = W0_addr[25:0];
  assign mem_130_4_W0_clk = W0_clk;
  assign mem_130_4_W0_data = W0_data[39:32];
  assign mem_130_4_W0_en = W0_en & W0_addr_sel == 8'h82;
  assign mem_130_4_W0_mask = W0_mask[4];
  assign mem_130_5_R0_addr = R0_addr[25:0];
  assign mem_130_5_R0_clk = R0_clk;
  assign mem_130_5_R0_en = R0_en & R0_addr_sel == 8'h82;
  assign mem_130_5_W0_addr = W0_addr[25:0];
  assign mem_130_5_W0_clk = W0_clk;
  assign mem_130_5_W0_data = W0_data[47:40];
  assign mem_130_5_W0_en = W0_en & W0_addr_sel == 8'h82;
  assign mem_130_5_W0_mask = W0_mask[5];
  assign mem_130_6_R0_addr = R0_addr[25:0];
  assign mem_130_6_R0_clk = R0_clk;
  assign mem_130_6_R0_en = R0_en & R0_addr_sel == 8'h82;
  assign mem_130_6_W0_addr = W0_addr[25:0];
  assign mem_130_6_W0_clk = W0_clk;
  assign mem_130_6_W0_data = W0_data[55:48];
  assign mem_130_6_W0_en = W0_en & W0_addr_sel == 8'h82;
  assign mem_130_6_W0_mask = W0_mask[6];
  assign mem_130_7_R0_addr = R0_addr[25:0];
  assign mem_130_7_R0_clk = R0_clk;
  assign mem_130_7_R0_en = R0_en & R0_addr_sel == 8'h82;
  assign mem_130_7_W0_addr = W0_addr[25:0];
  assign mem_130_7_W0_clk = W0_clk;
  assign mem_130_7_W0_data = W0_data[63:56];
  assign mem_130_7_W0_en = W0_en & W0_addr_sel == 8'h82;
  assign mem_130_7_W0_mask = W0_mask[7];
  assign mem_131_0_R0_addr = R0_addr[25:0];
  assign mem_131_0_R0_clk = R0_clk;
  assign mem_131_0_R0_en = R0_en & R0_addr_sel == 8'h83;
  assign mem_131_0_W0_addr = W0_addr[25:0];
  assign mem_131_0_W0_clk = W0_clk;
  assign mem_131_0_W0_data = W0_data[7:0];
  assign mem_131_0_W0_en = W0_en & W0_addr_sel == 8'h83;
  assign mem_131_0_W0_mask = W0_mask[0];
  assign mem_131_1_R0_addr = R0_addr[25:0];
  assign mem_131_1_R0_clk = R0_clk;
  assign mem_131_1_R0_en = R0_en & R0_addr_sel == 8'h83;
  assign mem_131_1_W0_addr = W0_addr[25:0];
  assign mem_131_1_W0_clk = W0_clk;
  assign mem_131_1_W0_data = W0_data[15:8];
  assign mem_131_1_W0_en = W0_en & W0_addr_sel == 8'h83;
  assign mem_131_1_W0_mask = W0_mask[1];
  assign mem_131_2_R0_addr = R0_addr[25:0];
  assign mem_131_2_R0_clk = R0_clk;
  assign mem_131_2_R0_en = R0_en & R0_addr_sel == 8'h83;
  assign mem_131_2_W0_addr = W0_addr[25:0];
  assign mem_131_2_W0_clk = W0_clk;
  assign mem_131_2_W0_data = W0_data[23:16];
  assign mem_131_2_W0_en = W0_en & W0_addr_sel == 8'h83;
  assign mem_131_2_W0_mask = W0_mask[2];
  assign mem_131_3_R0_addr = R0_addr[25:0];
  assign mem_131_3_R0_clk = R0_clk;
  assign mem_131_3_R0_en = R0_en & R0_addr_sel == 8'h83;
  assign mem_131_3_W0_addr = W0_addr[25:0];
  assign mem_131_3_W0_clk = W0_clk;
  assign mem_131_3_W0_data = W0_data[31:24];
  assign mem_131_3_W0_en = W0_en & W0_addr_sel == 8'h83;
  assign mem_131_3_W0_mask = W0_mask[3];
  assign mem_131_4_R0_addr = R0_addr[25:0];
  assign mem_131_4_R0_clk = R0_clk;
  assign mem_131_4_R0_en = R0_en & R0_addr_sel == 8'h83;
  assign mem_131_4_W0_addr = W0_addr[25:0];
  assign mem_131_4_W0_clk = W0_clk;
  assign mem_131_4_W0_data = W0_data[39:32];
  assign mem_131_4_W0_en = W0_en & W0_addr_sel == 8'h83;
  assign mem_131_4_W0_mask = W0_mask[4];
  assign mem_131_5_R0_addr = R0_addr[25:0];
  assign mem_131_5_R0_clk = R0_clk;
  assign mem_131_5_R0_en = R0_en & R0_addr_sel == 8'h83;
  assign mem_131_5_W0_addr = W0_addr[25:0];
  assign mem_131_5_W0_clk = W0_clk;
  assign mem_131_5_W0_data = W0_data[47:40];
  assign mem_131_5_W0_en = W0_en & W0_addr_sel == 8'h83;
  assign mem_131_5_W0_mask = W0_mask[5];
  assign mem_131_6_R0_addr = R0_addr[25:0];
  assign mem_131_6_R0_clk = R0_clk;
  assign mem_131_6_R0_en = R0_en & R0_addr_sel == 8'h83;
  assign mem_131_6_W0_addr = W0_addr[25:0];
  assign mem_131_6_W0_clk = W0_clk;
  assign mem_131_6_W0_data = W0_data[55:48];
  assign mem_131_6_W0_en = W0_en & W0_addr_sel == 8'h83;
  assign mem_131_6_W0_mask = W0_mask[6];
  assign mem_131_7_R0_addr = R0_addr[25:0];
  assign mem_131_7_R0_clk = R0_clk;
  assign mem_131_7_R0_en = R0_en & R0_addr_sel == 8'h83;
  assign mem_131_7_W0_addr = W0_addr[25:0];
  assign mem_131_7_W0_clk = W0_clk;
  assign mem_131_7_W0_data = W0_data[63:56];
  assign mem_131_7_W0_en = W0_en & W0_addr_sel == 8'h83;
  assign mem_131_7_W0_mask = W0_mask[7];
  assign mem_132_0_R0_addr = R0_addr[25:0];
  assign mem_132_0_R0_clk = R0_clk;
  assign mem_132_0_R0_en = R0_en & R0_addr_sel == 8'h84;
  assign mem_132_0_W0_addr = W0_addr[25:0];
  assign mem_132_0_W0_clk = W0_clk;
  assign mem_132_0_W0_data = W0_data[7:0];
  assign mem_132_0_W0_en = W0_en & W0_addr_sel == 8'h84;
  assign mem_132_0_W0_mask = W0_mask[0];
  assign mem_132_1_R0_addr = R0_addr[25:0];
  assign mem_132_1_R0_clk = R0_clk;
  assign mem_132_1_R0_en = R0_en & R0_addr_sel == 8'h84;
  assign mem_132_1_W0_addr = W0_addr[25:0];
  assign mem_132_1_W0_clk = W0_clk;
  assign mem_132_1_W0_data = W0_data[15:8];
  assign mem_132_1_W0_en = W0_en & W0_addr_sel == 8'h84;
  assign mem_132_1_W0_mask = W0_mask[1];
  assign mem_132_2_R0_addr = R0_addr[25:0];
  assign mem_132_2_R0_clk = R0_clk;
  assign mem_132_2_R0_en = R0_en & R0_addr_sel == 8'h84;
  assign mem_132_2_W0_addr = W0_addr[25:0];
  assign mem_132_2_W0_clk = W0_clk;
  assign mem_132_2_W0_data = W0_data[23:16];
  assign mem_132_2_W0_en = W0_en & W0_addr_sel == 8'h84;
  assign mem_132_2_W0_mask = W0_mask[2];
  assign mem_132_3_R0_addr = R0_addr[25:0];
  assign mem_132_3_R0_clk = R0_clk;
  assign mem_132_3_R0_en = R0_en & R0_addr_sel == 8'h84;
  assign mem_132_3_W0_addr = W0_addr[25:0];
  assign mem_132_3_W0_clk = W0_clk;
  assign mem_132_3_W0_data = W0_data[31:24];
  assign mem_132_3_W0_en = W0_en & W0_addr_sel == 8'h84;
  assign mem_132_3_W0_mask = W0_mask[3];
  assign mem_132_4_R0_addr = R0_addr[25:0];
  assign mem_132_4_R0_clk = R0_clk;
  assign mem_132_4_R0_en = R0_en & R0_addr_sel == 8'h84;
  assign mem_132_4_W0_addr = W0_addr[25:0];
  assign mem_132_4_W0_clk = W0_clk;
  assign mem_132_4_W0_data = W0_data[39:32];
  assign mem_132_4_W0_en = W0_en & W0_addr_sel == 8'h84;
  assign mem_132_4_W0_mask = W0_mask[4];
  assign mem_132_5_R0_addr = R0_addr[25:0];
  assign mem_132_5_R0_clk = R0_clk;
  assign mem_132_5_R0_en = R0_en & R0_addr_sel == 8'h84;
  assign mem_132_5_W0_addr = W0_addr[25:0];
  assign mem_132_5_W0_clk = W0_clk;
  assign mem_132_5_W0_data = W0_data[47:40];
  assign mem_132_5_W0_en = W0_en & W0_addr_sel == 8'h84;
  assign mem_132_5_W0_mask = W0_mask[5];
  assign mem_132_6_R0_addr = R0_addr[25:0];
  assign mem_132_6_R0_clk = R0_clk;
  assign mem_132_6_R0_en = R0_en & R0_addr_sel == 8'h84;
  assign mem_132_6_W0_addr = W0_addr[25:0];
  assign mem_132_6_W0_clk = W0_clk;
  assign mem_132_6_W0_data = W0_data[55:48];
  assign mem_132_6_W0_en = W0_en & W0_addr_sel == 8'h84;
  assign mem_132_6_W0_mask = W0_mask[6];
  assign mem_132_7_R0_addr = R0_addr[25:0];
  assign mem_132_7_R0_clk = R0_clk;
  assign mem_132_7_R0_en = R0_en & R0_addr_sel == 8'h84;
  assign mem_132_7_W0_addr = W0_addr[25:0];
  assign mem_132_7_W0_clk = W0_clk;
  assign mem_132_7_W0_data = W0_data[63:56];
  assign mem_132_7_W0_en = W0_en & W0_addr_sel == 8'h84;
  assign mem_132_7_W0_mask = W0_mask[7];
  assign mem_133_0_R0_addr = R0_addr[25:0];
  assign mem_133_0_R0_clk = R0_clk;
  assign mem_133_0_R0_en = R0_en & R0_addr_sel == 8'h85;
  assign mem_133_0_W0_addr = W0_addr[25:0];
  assign mem_133_0_W0_clk = W0_clk;
  assign mem_133_0_W0_data = W0_data[7:0];
  assign mem_133_0_W0_en = W0_en & W0_addr_sel == 8'h85;
  assign mem_133_0_W0_mask = W0_mask[0];
  assign mem_133_1_R0_addr = R0_addr[25:0];
  assign mem_133_1_R0_clk = R0_clk;
  assign mem_133_1_R0_en = R0_en & R0_addr_sel == 8'h85;
  assign mem_133_1_W0_addr = W0_addr[25:0];
  assign mem_133_1_W0_clk = W0_clk;
  assign mem_133_1_W0_data = W0_data[15:8];
  assign mem_133_1_W0_en = W0_en & W0_addr_sel == 8'h85;
  assign mem_133_1_W0_mask = W0_mask[1];
  assign mem_133_2_R0_addr = R0_addr[25:0];
  assign mem_133_2_R0_clk = R0_clk;
  assign mem_133_2_R0_en = R0_en & R0_addr_sel == 8'h85;
  assign mem_133_2_W0_addr = W0_addr[25:0];
  assign mem_133_2_W0_clk = W0_clk;
  assign mem_133_2_W0_data = W0_data[23:16];
  assign mem_133_2_W0_en = W0_en & W0_addr_sel == 8'h85;
  assign mem_133_2_W0_mask = W0_mask[2];
  assign mem_133_3_R0_addr = R0_addr[25:0];
  assign mem_133_3_R0_clk = R0_clk;
  assign mem_133_3_R0_en = R0_en & R0_addr_sel == 8'h85;
  assign mem_133_3_W0_addr = W0_addr[25:0];
  assign mem_133_3_W0_clk = W0_clk;
  assign mem_133_3_W0_data = W0_data[31:24];
  assign mem_133_3_W0_en = W0_en & W0_addr_sel == 8'h85;
  assign mem_133_3_W0_mask = W0_mask[3];
  assign mem_133_4_R0_addr = R0_addr[25:0];
  assign mem_133_4_R0_clk = R0_clk;
  assign mem_133_4_R0_en = R0_en & R0_addr_sel == 8'h85;
  assign mem_133_4_W0_addr = W0_addr[25:0];
  assign mem_133_4_W0_clk = W0_clk;
  assign mem_133_4_W0_data = W0_data[39:32];
  assign mem_133_4_W0_en = W0_en & W0_addr_sel == 8'h85;
  assign mem_133_4_W0_mask = W0_mask[4];
  assign mem_133_5_R0_addr = R0_addr[25:0];
  assign mem_133_5_R0_clk = R0_clk;
  assign mem_133_5_R0_en = R0_en & R0_addr_sel == 8'h85;
  assign mem_133_5_W0_addr = W0_addr[25:0];
  assign mem_133_5_W0_clk = W0_clk;
  assign mem_133_5_W0_data = W0_data[47:40];
  assign mem_133_5_W0_en = W0_en & W0_addr_sel == 8'h85;
  assign mem_133_5_W0_mask = W0_mask[5];
  assign mem_133_6_R0_addr = R0_addr[25:0];
  assign mem_133_6_R0_clk = R0_clk;
  assign mem_133_6_R0_en = R0_en & R0_addr_sel == 8'h85;
  assign mem_133_6_W0_addr = W0_addr[25:0];
  assign mem_133_6_W0_clk = W0_clk;
  assign mem_133_6_W0_data = W0_data[55:48];
  assign mem_133_6_W0_en = W0_en & W0_addr_sel == 8'h85;
  assign mem_133_6_W0_mask = W0_mask[6];
  assign mem_133_7_R0_addr = R0_addr[25:0];
  assign mem_133_7_R0_clk = R0_clk;
  assign mem_133_7_R0_en = R0_en & R0_addr_sel == 8'h85;
  assign mem_133_7_W0_addr = W0_addr[25:0];
  assign mem_133_7_W0_clk = W0_clk;
  assign mem_133_7_W0_data = W0_data[63:56];
  assign mem_133_7_W0_en = W0_en & W0_addr_sel == 8'h85;
  assign mem_133_7_W0_mask = W0_mask[7];
  assign mem_134_0_R0_addr = R0_addr[25:0];
  assign mem_134_0_R0_clk = R0_clk;
  assign mem_134_0_R0_en = R0_en & R0_addr_sel == 8'h86;
  assign mem_134_0_W0_addr = W0_addr[25:0];
  assign mem_134_0_W0_clk = W0_clk;
  assign mem_134_0_W0_data = W0_data[7:0];
  assign mem_134_0_W0_en = W0_en & W0_addr_sel == 8'h86;
  assign mem_134_0_W0_mask = W0_mask[0];
  assign mem_134_1_R0_addr = R0_addr[25:0];
  assign mem_134_1_R0_clk = R0_clk;
  assign mem_134_1_R0_en = R0_en & R0_addr_sel == 8'h86;
  assign mem_134_1_W0_addr = W0_addr[25:0];
  assign mem_134_1_W0_clk = W0_clk;
  assign mem_134_1_W0_data = W0_data[15:8];
  assign mem_134_1_W0_en = W0_en & W0_addr_sel == 8'h86;
  assign mem_134_1_W0_mask = W0_mask[1];
  assign mem_134_2_R0_addr = R0_addr[25:0];
  assign mem_134_2_R0_clk = R0_clk;
  assign mem_134_2_R0_en = R0_en & R0_addr_sel == 8'h86;
  assign mem_134_2_W0_addr = W0_addr[25:0];
  assign mem_134_2_W0_clk = W0_clk;
  assign mem_134_2_W0_data = W0_data[23:16];
  assign mem_134_2_W0_en = W0_en & W0_addr_sel == 8'h86;
  assign mem_134_2_W0_mask = W0_mask[2];
  assign mem_134_3_R0_addr = R0_addr[25:0];
  assign mem_134_3_R0_clk = R0_clk;
  assign mem_134_3_R0_en = R0_en & R0_addr_sel == 8'h86;
  assign mem_134_3_W0_addr = W0_addr[25:0];
  assign mem_134_3_W0_clk = W0_clk;
  assign mem_134_3_W0_data = W0_data[31:24];
  assign mem_134_3_W0_en = W0_en & W0_addr_sel == 8'h86;
  assign mem_134_3_W0_mask = W0_mask[3];
  assign mem_134_4_R0_addr = R0_addr[25:0];
  assign mem_134_4_R0_clk = R0_clk;
  assign mem_134_4_R0_en = R0_en & R0_addr_sel == 8'h86;
  assign mem_134_4_W0_addr = W0_addr[25:0];
  assign mem_134_4_W0_clk = W0_clk;
  assign mem_134_4_W0_data = W0_data[39:32];
  assign mem_134_4_W0_en = W0_en & W0_addr_sel == 8'h86;
  assign mem_134_4_W0_mask = W0_mask[4];
  assign mem_134_5_R0_addr = R0_addr[25:0];
  assign mem_134_5_R0_clk = R0_clk;
  assign mem_134_5_R0_en = R0_en & R0_addr_sel == 8'h86;
  assign mem_134_5_W0_addr = W0_addr[25:0];
  assign mem_134_5_W0_clk = W0_clk;
  assign mem_134_5_W0_data = W0_data[47:40];
  assign mem_134_5_W0_en = W0_en & W0_addr_sel == 8'h86;
  assign mem_134_5_W0_mask = W0_mask[5];
  assign mem_134_6_R0_addr = R0_addr[25:0];
  assign mem_134_6_R0_clk = R0_clk;
  assign mem_134_6_R0_en = R0_en & R0_addr_sel == 8'h86;
  assign mem_134_6_W0_addr = W0_addr[25:0];
  assign mem_134_6_W0_clk = W0_clk;
  assign mem_134_6_W0_data = W0_data[55:48];
  assign mem_134_6_W0_en = W0_en & W0_addr_sel == 8'h86;
  assign mem_134_6_W0_mask = W0_mask[6];
  assign mem_134_7_R0_addr = R0_addr[25:0];
  assign mem_134_7_R0_clk = R0_clk;
  assign mem_134_7_R0_en = R0_en & R0_addr_sel == 8'h86;
  assign mem_134_7_W0_addr = W0_addr[25:0];
  assign mem_134_7_W0_clk = W0_clk;
  assign mem_134_7_W0_data = W0_data[63:56];
  assign mem_134_7_W0_en = W0_en & W0_addr_sel == 8'h86;
  assign mem_134_7_W0_mask = W0_mask[7];
  assign mem_135_0_R0_addr = R0_addr[25:0];
  assign mem_135_0_R0_clk = R0_clk;
  assign mem_135_0_R0_en = R0_en & R0_addr_sel == 8'h87;
  assign mem_135_0_W0_addr = W0_addr[25:0];
  assign mem_135_0_W0_clk = W0_clk;
  assign mem_135_0_W0_data = W0_data[7:0];
  assign mem_135_0_W0_en = W0_en & W0_addr_sel == 8'h87;
  assign mem_135_0_W0_mask = W0_mask[0];
  assign mem_135_1_R0_addr = R0_addr[25:0];
  assign mem_135_1_R0_clk = R0_clk;
  assign mem_135_1_R0_en = R0_en & R0_addr_sel == 8'h87;
  assign mem_135_1_W0_addr = W0_addr[25:0];
  assign mem_135_1_W0_clk = W0_clk;
  assign mem_135_1_W0_data = W0_data[15:8];
  assign mem_135_1_W0_en = W0_en & W0_addr_sel == 8'h87;
  assign mem_135_1_W0_mask = W0_mask[1];
  assign mem_135_2_R0_addr = R0_addr[25:0];
  assign mem_135_2_R0_clk = R0_clk;
  assign mem_135_2_R0_en = R0_en & R0_addr_sel == 8'h87;
  assign mem_135_2_W0_addr = W0_addr[25:0];
  assign mem_135_2_W0_clk = W0_clk;
  assign mem_135_2_W0_data = W0_data[23:16];
  assign mem_135_2_W0_en = W0_en & W0_addr_sel == 8'h87;
  assign mem_135_2_W0_mask = W0_mask[2];
  assign mem_135_3_R0_addr = R0_addr[25:0];
  assign mem_135_3_R0_clk = R0_clk;
  assign mem_135_3_R0_en = R0_en & R0_addr_sel == 8'h87;
  assign mem_135_3_W0_addr = W0_addr[25:0];
  assign mem_135_3_W0_clk = W0_clk;
  assign mem_135_3_W0_data = W0_data[31:24];
  assign mem_135_3_W0_en = W0_en & W0_addr_sel == 8'h87;
  assign mem_135_3_W0_mask = W0_mask[3];
  assign mem_135_4_R0_addr = R0_addr[25:0];
  assign mem_135_4_R0_clk = R0_clk;
  assign mem_135_4_R0_en = R0_en & R0_addr_sel == 8'h87;
  assign mem_135_4_W0_addr = W0_addr[25:0];
  assign mem_135_4_W0_clk = W0_clk;
  assign mem_135_4_W0_data = W0_data[39:32];
  assign mem_135_4_W0_en = W0_en & W0_addr_sel == 8'h87;
  assign mem_135_4_W0_mask = W0_mask[4];
  assign mem_135_5_R0_addr = R0_addr[25:0];
  assign mem_135_5_R0_clk = R0_clk;
  assign mem_135_5_R0_en = R0_en & R0_addr_sel == 8'h87;
  assign mem_135_5_W0_addr = W0_addr[25:0];
  assign mem_135_5_W0_clk = W0_clk;
  assign mem_135_5_W0_data = W0_data[47:40];
  assign mem_135_5_W0_en = W0_en & W0_addr_sel == 8'h87;
  assign mem_135_5_W0_mask = W0_mask[5];
  assign mem_135_6_R0_addr = R0_addr[25:0];
  assign mem_135_6_R0_clk = R0_clk;
  assign mem_135_6_R0_en = R0_en & R0_addr_sel == 8'h87;
  assign mem_135_6_W0_addr = W0_addr[25:0];
  assign mem_135_6_W0_clk = W0_clk;
  assign mem_135_6_W0_data = W0_data[55:48];
  assign mem_135_6_W0_en = W0_en & W0_addr_sel == 8'h87;
  assign mem_135_6_W0_mask = W0_mask[6];
  assign mem_135_7_R0_addr = R0_addr[25:0];
  assign mem_135_7_R0_clk = R0_clk;
  assign mem_135_7_R0_en = R0_en & R0_addr_sel == 8'h87;
  assign mem_135_7_W0_addr = W0_addr[25:0];
  assign mem_135_7_W0_clk = W0_clk;
  assign mem_135_7_W0_data = W0_data[63:56];
  assign mem_135_7_W0_en = W0_en & W0_addr_sel == 8'h87;
  assign mem_135_7_W0_mask = W0_mask[7];
  assign mem_136_0_R0_addr = R0_addr[25:0];
  assign mem_136_0_R0_clk = R0_clk;
  assign mem_136_0_R0_en = R0_en & R0_addr_sel == 8'h88;
  assign mem_136_0_W0_addr = W0_addr[25:0];
  assign mem_136_0_W0_clk = W0_clk;
  assign mem_136_0_W0_data = W0_data[7:0];
  assign mem_136_0_W0_en = W0_en & W0_addr_sel == 8'h88;
  assign mem_136_0_W0_mask = W0_mask[0];
  assign mem_136_1_R0_addr = R0_addr[25:0];
  assign mem_136_1_R0_clk = R0_clk;
  assign mem_136_1_R0_en = R0_en & R0_addr_sel == 8'h88;
  assign mem_136_1_W0_addr = W0_addr[25:0];
  assign mem_136_1_W0_clk = W0_clk;
  assign mem_136_1_W0_data = W0_data[15:8];
  assign mem_136_1_W0_en = W0_en & W0_addr_sel == 8'h88;
  assign mem_136_1_W0_mask = W0_mask[1];
  assign mem_136_2_R0_addr = R0_addr[25:0];
  assign mem_136_2_R0_clk = R0_clk;
  assign mem_136_2_R0_en = R0_en & R0_addr_sel == 8'h88;
  assign mem_136_2_W0_addr = W0_addr[25:0];
  assign mem_136_2_W0_clk = W0_clk;
  assign mem_136_2_W0_data = W0_data[23:16];
  assign mem_136_2_W0_en = W0_en & W0_addr_sel == 8'h88;
  assign mem_136_2_W0_mask = W0_mask[2];
  assign mem_136_3_R0_addr = R0_addr[25:0];
  assign mem_136_3_R0_clk = R0_clk;
  assign mem_136_3_R0_en = R0_en & R0_addr_sel == 8'h88;
  assign mem_136_3_W0_addr = W0_addr[25:0];
  assign mem_136_3_W0_clk = W0_clk;
  assign mem_136_3_W0_data = W0_data[31:24];
  assign mem_136_3_W0_en = W0_en & W0_addr_sel == 8'h88;
  assign mem_136_3_W0_mask = W0_mask[3];
  assign mem_136_4_R0_addr = R0_addr[25:0];
  assign mem_136_4_R0_clk = R0_clk;
  assign mem_136_4_R0_en = R0_en & R0_addr_sel == 8'h88;
  assign mem_136_4_W0_addr = W0_addr[25:0];
  assign mem_136_4_W0_clk = W0_clk;
  assign mem_136_4_W0_data = W0_data[39:32];
  assign mem_136_4_W0_en = W0_en & W0_addr_sel == 8'h88;
  assign mem_136_4_W0_mask = W0_mask[4];
  assign mem_136_5_R0_addr = R0_addr[25:0];
  assign mem_136_5_R0_clk = R0_clk;
  assign mem_136_5_R0_en = R0_en & R0_addr_sel == 8'h88;
  assign mem_136_5_W0_addr = W0_addr[25:0];
  assign mem_136_5_W0_clk = W0_clk;
  assign mem_136_5_W0_data = W0_data[47:40];
  assign mem_136_5_W0_en = W0_en & W0_addr_sel == 8'h88;
  assign mem_136_5_W0_mask = W0_mask[5];
  assign mem_136_6_R0_addr = R0_addr[25:0];
  assign mem_136_6_R0_clk = R0_clk;
  assign mem_136_6_R0_en = R0_en & R0_addr_sel == 8'h88;
  assign mem_136_6_W0_addr = W0_addr[25:0];
  assign mem_136_6_W0_clk = W0_clk;
  assign mem_136_6_W0_data = W0_data[55:48];
  assign mem_136_6_W0_en = W0_en & W0_addr_sel == 8'h88;
  assign mem_136_6_W0_mask = W0_mask[6];
  assign mem_136_7_R0_addr = R0_addr[25:0];
  assign mem_136_7_R0_clk = R0_clk;
  assign mem_136_7_R0_en = R0_en & R0_addr_sel == 8'h88;
  assign mem_136_7_W0_addr = W0_addr[25:0];
  assign mem_136_7_W0_clk = W0_clk;
  assign mem_136_7_W0_data = W0_data[63:56];
  assign mem_136_7_W0_en = W0_en & W0_addr_sel == 8'h88;
  assign mem_136_7_W0_mask = W0_mask[7];
  assign mem_137_0_R0_addr = R0_addr[25:0];
  assign mem_137_0_R0_clk = R0_clk;
  assign mem_137_0_R0_en = R0_en & R0_addr_sel == 8'h89;
  assign mem_137_0_W0_addr = W0_addr[25:0];
  assign mem_137_0_W0_clk = W0_clk;
  assign mem_137_0_W0_data = W0_data[7:0];
  assign mem_137_0_W0_en = W0_en & W0_addr_sel == 8'h89;
  assign mem_137_0_W0_mask = W0_mask[0];
  assign mem_137_1_R0_addr = R0_addr[25:0];
  assign mem_137_1_R0_clk = R0_clk;
  assign mem_137_1_R0_en = R0_en & R0_addr_sel == 8'h89;
  assign mem_137_1_W0_addr = W0_addr[25:0];
  assign mem_137_1_W0_clk = W0_clk;
  assign mem_137_1_W0_data = W0_data[15:8];
  assign mem_137_1_W0_en = W0_en & W0_addr_sel == 8'h89;
  assign mem_137_1_W0_mask = W0_mask[1];
  assign mem_137_2_R0_addr = R0_addr[25:0];
  assign mem_137_2_R0_clk = R0_clk;
  assign mem_137_2_R0_en = R0_en & R0_addr_sel == 8'h89;
  assign mem_137_2_W0_addr = W0_addr[25:0];
  assign mem_137_2_W0_clk = W0_clk;
  assign mem_137_2_W0_data = W0_data[23:16];
  assign mem_137_2_W0_en = W0_en & W0_addr_sel == 8'h89;
  assign mem_137_2_W0_mask = W0_mask[2];
  assign mem_137_3_R0_addr = R0_addr[25:0];
  assign mem_137_3_R0_clk = R0_clk;
  assign mem_137_3_R0_en = R0_en & R0_addr_sel == 8'h89;
  assign mem_137_3_W0_addr = W0_addr[25:0];
  assign mem_137_3_W0_clk = W0_clk;
  assign mem_137_3_W0_data = W0_data[31:24];
  assign mem_137_3_W0_en = W0_en & W0_addr_sel == 8'h89;
  assign mem_137_3_W0_mask = W0_mask[3];
  assign mem_137_4_R0_addr = R0_addr[25:0];
  assign mem_137_4_R0_clk = R0_clk;
  assign mem_137_4_R0_en = R0_en & R0_addr_sel == 8'h89;
  assign mem_137_4_W0_addr = W0_addr[25:0];
  assign mem_137_4_W0_clk = W0_clk;
  assign mem_137_4_W0_data = W0_data[39:32];
  assign mem_137_4_W0_en = W0_en & W0_addr_sel == 8'h89;
  assign mem_137_4_W0_mask = W0_mask[4];
  assign mem_137_5_R0_addr = R0_addr[25:0];
  assign mem_137_5_R0_clk = R0_clk;
  assign mem_137_5_R0_en = R0_en & R0_addr_sel == 8'h89;
  assign mem_137_5_W0_addr = W0_addr[25:0];
  assign mem_137_5_W0_clk = W0_clk;
  assign mem_137_5_W0_data = W0_data[47:40];
  assign mem_137_5_W0_en = W0_en & W0_addr_sel == 8'h89;
  assign mem_137_5_W0_mask = W0_mask[5];
  assign mem_137_6_R0_addr = R0_addr[25:0];
  assign mem_137_6_R0_clk = R0_clk;
  assign mem_137_6_R0_en = R0_en & R0_addr_sel == 8'h89;
  assign mem_137_6_W0_addr = W0_addr[25:0];
  assign mem_137_6_W0_clk = W0_clk;
  assign mem_137_6_W0_data = W0_data[55:48];
  assign mem_137_6_W0_en = W0_en & W0_addr_sel == 8'h89;
  assign mem_137_6_W0_mask = W0_mask[6];
  assign mem_137_7_R0_addr = R0_addr[25:0];
  assign mem_137_7_R0_clk = R0_clk;
  assign mem_137_7_R0_en = R0_en & R0_addr_sel == 8'h89;
  assign mem_137_7_W0_addr = W0_addr[25:0];
  assign mem_137_7_W0_clk = W0_clk;
  assign mem_137_7_W0_data = W0_data[63:56];
  assign mem_137_7_W0_en = W0_en & W0_addr_sel == 8'h89;
  assign mem_137_7_W0_mask = W0_mask[7];
  assign mem_138_0_R0_addr = R0_addr[25:0];
  assign mem_138_0_R0_clk = R0_clk;
  assign mem_138_0_R0_en = R0_en & R0_addr_sel == 8'h8a;
  assign mem_138_0_W0_addr = W0_addr[25:0];
  assign mem_138_0_W0_clk = W0_clk;
  assign mem_138_0_W0_data = W0_data[7:0];
  assign mem_138_0_W0_en = W0_en & W0_addr_sel == 8'h8a;
  assign mem_138_0_W0_mask = W0_mask[0];
  assign mem_138_1_R0_addr = R0_addr[25:0];
  assign mem_138_1_R0_clk = R0_clk;
  assign mem_138_1_R0_en = R0_en & R0_addr_sel == 8'h8a;
  assign mem_138_1_W0_addr = W0_addr[25:0];
  assign mem_138_1_W0_clk = W0_clk;
  assign mem_138_1_W0_data = W0_data[15:8];
  assign mem_138_1_W0_en = W0_en & W0_addr_sel == 8'h8a;
  assign mem_138_1_W0_mask = W0_mask[1];
  assign mem_138_2_R0_addr = R0_addr[25:0];
  assign mem_138_2_R0_clk = R0_clk;
  assign mem_138_2_R0_en = R0_en & R0_addr_sel == 8'h8a;
  assign mem_138_2_W0_addr = W0_addr[25:0];
  assign mem_138_2_W0_clk = W0_clk;
  assign mem_138_2_W0_data = W0_data[23:16];
  assign mem_138_2_W0_en = W0_en & W0_addr_sel == 8'h8a;
  assign mem_138_2_W0_mask = W0_mask[2];
  assign mem_138_3_R0_addr = R0_addr[25:0];
  assign mem_138_3_R0_clk = R0_clk;
  assign mem_138_3_R0_en = R0_en & R0_addr_sel == 8'h8a;
  assign mem_138_3_W0_addr = W0_addr[25:0];
  assign mem_138_3_W0_clk = W0_clk;
  assign mem_138_3_W0_data = W0_data[31:24];
  assign mem_138_3_W0_en = W0_en & W0_addr_sel == 8'h8a;
  assign mem_138_3_W0_mask = W0_mask[3];
  assign mem_138_4_R0_addr = R0_addr[25:0];
  assign mem_138_4_R0_clk = R0_clk;
  assign mem_138_4_R0_en = R0_en & R0_addr_sel == 8'h8a;
  assign mem_138_4_W0_addr = W0_addr[25:0];
  assign mem_138_4_W0_clk = W0_clk;
  assign mem_138_4_W0_data = W0_data[39:32];
  assign mem_138_4_W0_en = W0_en & W0_addr_sel == 8'h8a;
  assign mem_138_4_W0_mask = W0_mask[4];
  assign mem_138_5_R0_addr = R0_addr[25:0];
  assign mem_138_5_R0_clk = R0_clk;
  assign mem_138_5_R0_en = R0_en & R0_addr_sel == 8'h8a;
  assign mem_138_5_W0_addr = W0_addr[25:0];
  assign mem_138_5_W0_clk = W0_clk;
  assign mem_138_5_W0_data = W0_data[47:40];
  assign mem_138_5_W0_en = W0_en & W0_addr_sel == 8'h8a;
  assign mem_138_5_W0_mask = W0_mask[5];
  assign mem_138_6_R0_addr = R0_addr[25:0];
  assign mem_138_6_R0_clk = R0_clk;
  assign mem_138_6_R0_en = R0_en & R0_addr_sel == 8'h8a;
  assign mem_138_6_W0_addr = W0_addr[25:0];
  assign mem_138_6_W0_clk = W0_clk;
  assign mem_138_6_W0_data = W0_data[55:48];
  assign mem_138_6_W0_en = W0_en & W0_addr_sel == 8'h8a;
  assign mem_138_6_W0_mask = W0_mask[6];
  assign mem_138_7_R0_addr = R0_addr[25:0];
  assign mem_138_7_R0_clk = R0_clk;
  assign mem_138_7_R0_en = R0_en & R0_addr_sel == 8'h8a;
  assign mem_138_7_W0_addr = W0_addr[25:0];
  assign mem_138_7_W0_clk = W0_clk;
  assign mem_138_7_W0_data = W0_data[63:56];
  assign mem_138_7_W0_en = W0_en & W0_addr_sel == 8'h8a;
  assign mem_138_7_W0_mask = W0_mask[7];
  assign mem_139_0_R0_addr = R0_addr[25:0];
  assign mem_139_0_R0_clk = R0_clk;
  assign mem_139_0_R0_en = R0_en & R0_addr_sel == 8'h8b;
  assign mem_139_0_W0_addr = W0_addr[25:0];
  assign mem_139_0_W0_clk = W0_clk;
  assign mem_139_0_W0_data = W0_data[7:0];
  assign mem_139_0_W0_en = W0_en & W0_addr_sel == 8'h8b;
  assign mem_139_0_W0_mask = W0_mask[0];
  assign mem_139_1_R0_addr = R0_addr[25:0];
  assign mem_139_1_R0_clk = R0_clk;
  assign mem_139_1_R0_en = R0_en & R0_addr_sel == 8'h8b;
  assign mem_139_1_W0_addr = W0_addr[25:0];
  assign mem_139_1_W0_clk = W0_clk;
  assign mem_139_1_W0_data = W0_data[15:8];
  assign mem_139_1_W0_en = W0_en & W0_addr_sel == 8'h8b;
  assign mem_139_1_W0_mask = W0_mask[1];
  assign mem_139_2_R0_addr = R0_addr[25:0];
  assign mem_139_2_R0_clk = R0_clk;
  assign mem_139_2_R0_en = R0_en & R0_addr_sel == 8'h8b;
  assign mem_139_2_W0_addr = W0_addr[25:0];
  assign mem_139_2_W0_clk = W0_clk;
  assign mem_139_2_W0_data = W0_data[23:16];
  assign mem_139_2_W0_en = W0_en & W0_addr_sel == 8'h8b;
  assign mem_139_2_W0_mask = W0_mask[2];
  assign mem_139_3_R0_addr = R0_addr[25:0];
  assign mem_139_3_R0_clk = R0_clk;
  assign mem_139_3_R0_en = R0_en & R0_addr_sel == 8'h8b;
  assign mem_139_3_W0_addr = W0_addr[25:0];
  assign mem_139_3_W0_clk = W0_clk;
  assign mem_139_3_W0_data = W0_data[31:24];
  assign mem_139_3_W0_en = W0_en & W0_addr_sel == 8'h8b;
  assign mem_139_3_W0_mask = W0_mask[3];
  assign mem_139_4_R0_addr = R0_addr[25:0];
  assign mem_139_4_R0_clk = R0_clk;
  assign mem_139_4_R0_en = R0_en & R0_addr_sel == 8'h8b;
  assign mem_139_4_W0_addr = W0_addr[25:0];
  assign mem_139_4_W0_clk = W0_clk;
  assign mem_139_4_W0_data = W0_data[39:32];
  assign mem_139_4_W0_en = W0_en & W0_addr_sel == 8'h8b;
  assign mem_139_4_W0_mask = W0_mask[4];
  assign mem_139_5_R0_addr = R0_addr[25:0];
  assign mem_139_5_R0_clk = R0_clk;
  assign mem_139_5_R0_en = R0_en & R0_addr_sel == 8'h8b;
  assign mem_139_5_W0_addr = W0_addr[25:0];
  assign mem_139_5_W0_clk = W0_clk;
  assign mem_139_5_W0_data = W0_data[47:40];
  assign mem_139_5_W0_en = W0_en & W0_addr_sel == 8'h8b;
  assign mem_139_5_W0_mask = W0_mask[5];
  assign mem_139_6_R0_addr = R0_addr[25:0];
  assign mem_139_6_R0_clk = R0_clk;
  assign mem_139_6_R0_en = R0_en & R0_addr_sel == 8'h8b;
  assign mem_139_6_W0_addr = W0_addr[25:0];
  assign mem_139_6_W0_clk = W0_clk;
  assign mem_139_6_W0_data = W0_data[55:48];
  assign mem_139_6_W0_en = W0_en & W0_addr_sel == 8'h8b;
  assign mem_139_6_W0_mask = W0_mask[6];
  assign mem_139_7_R0_addr = R0_addr[25:0];
  assign mem_139_7_R0_clk = R0_clk;
  assign mem_139_7_R0_en = R0_en & R0_addr_sel == 8'h8b;
  assign mem_139_7_W0_addr = W0_addr[25:0];
  assign mem_139_7_W0_clk = W0_clk;
  assign mem_139_7_W0_data = W0_data[63:56];
  assign mem_139_7_W0_en = W0_en & W0_addr_sel == 8'h8b;
  assign mem_139_7_W0_mask = W0_mask[7];
  assign mem_140_0_R0_addr = R0_addr[25:0];
  assign mem_140_0_R0_clk = R0_clk;
  assign mem_140_0_R0_en = R0_en & R0_addr_sel == 8'h8c;
  assign mem_140_0_W0_addr = W0_addr[25:0];
  assign mem_140_0_W0_clk = W0_clk;
  assign mem_140_0_W0_data = W0_data[7:0];
  assign mem_140_0_W0_en = W0_en & W0_addr_sel == 8'h8c;
  assign mem_140_0_W0_mask = W0_mask[0];
  assign mem_140_1_R0_addr = R0_addr[25:0];
  assign mem_140_1_R0_clk = R0_clk;
  assign mem_140_1_R0_en = R0_en & R0_addr_sel == 8'h8c;
  assign mem_140_1_W0_addr = W0_addr[25:0];
  assign mem_140_1_W0_clk = W0_clk;
  assign mem_140_1_W0_data = W0_data[15:8];
  assign mem_140_1_W0_en = W0_en & W0_addr_sel == 8'h8c;
  assign mem_140_1_W0_mask = W0_mask[1];
  assign mem_140_2_R0_addr = R0_addr[25:0];
  assign mem_140_2_R0_clk = R0_clk;
  assign mem_140_2_R0_en = R0_en & R0_addr_sel == 8'h8c;
  assign mem_140_2_W0_addr = W0_addr[25:0];
  assign mem_140_2_W0_clk = W0_clk;
  assign mem_140_2_W0_data = W0_data[23:16];
  assign mem_140_2_W0_en = W0_en & W0_addr_sel == 8'h8c;
  assign mem_140_2_W0_mask = W0_mask[2];
  assign mem_140_3_R0_addr = R0_addr[25:0];
  assign mem_140_3_R0_clk = R0_clk;
  assign mem_140_3_R0_en = R0_en & R0_addr_sel == 8'h8c;
  assign mem_140_3_W0_addr = W0_addr[25:0];
  assign mem_140_3_W0_clk = W0_clk;
  assign mem_140_3_W0_data = W0_data[31:24];
  assign mem_140_3_W0_en = W0_en & W0_addr_sel == 8'h8c;
  assign mem_140_3_W0_mask = W0_mask[3];
  assign mem_140_4_R0_addr = R0_addr[25:0];
  assign mem_140_4_R0_clk = R0_clk;
  assign mem_140_4_R0_en = R0_en & R0_addr_sel == 8'h8c;
  assign mem_140_4_W0_addr = W0_addr[25:0];
  assign mem_140_4_W0_clk = W0_clk;
  assign mem_140_4_W0_data = W0_data[39:32];
  assign mem_140_4_W0_en = W0_en & W0_addr_sel == 8'h8c;
  assign mem_140_4_W0_mask = W0_mask[4];
  assign mem_140_5_R0_addr = R0_addr[25:0];
  assign mem_140_5_R0_clk = R0_clk;
  assign mem_140_5_R0_en = R0_en & R0_addr_sel == 8'h8c;
  assign mem_140_5_W0_addr = W0_addr[25:0];
  assign mem_140_5_W0_clk = W0_clk;
  assign mem_140_5_W0_data = W0_data[47:40];
  assign mem_140_5_W0_en = W0_en & W0_addr_sel == 8'h8c;
  assign mem_140_5_W0_mask = W0_mask[5];
  assign mem_140_6_R0_addr = R0_addr[25:0];
  assign mem_140_6_R0_clk = R0_clk;
  assign mem_140_6_R0_en = R0_en & R0_addr_sel == 8'h8c;
  assign mem_140_6_W0_addr = W0_addr[25:0];
  assign mem_140_6_W0_clk = W0_clk;
  assign mem_140_6_W0_data = W0_data[55:48];
  assign mem_140_6_W0_en = W0_en & W0_addr_sel == 8'h8c;
  assign mem_140_6_W0_mask = W0_mask[6];
  assign mem_140_7_R0_addr = R0_addr[25:0];
  assign mem_140_7_R0_clk = R0_clk;
  assign mem_140_7_R0_en = R0_en & R0_addr_sel == 8'h8c;
  assign mem_140_7_W0_addr = W0_addr[25:0];
  assign mem_140_7_W0_clk = W0_clk;
  assign mem_140_7_W0_data = W0_data[63:56];
  assign mem_140_7_W0_en = W0_en & W0_addr_sel == 8'h8c;
  assign mem_140_7_W0_mask = W0_mask[7];
  assign mem_141_0_R0_addr = R0_addr[25:0];
  assign mem_141_0_R0_clk = R0_clk;
  assign mem_141_0_R0_en = R0_en & R0_addr_sel == 8'h8d;
  assign mem_141_0_W0_addr = W0_addr[25:0];
  assign mem_141_0_W0_clk = W0_clk;
  assign mem_141_0_W0_data = W0_data[7:0];
  assign mem_141_0_W0_en = W0_en & W0_addr_sel == 8'h8d;
  assign mem_141_0_W0_mask = W0_mask[0];
  assign mem_141_1_R0_addr = R0_addr[25:0];
  assign mem_141_1_R0_clk = R0_clk;
  assign mem_141_1_R0_en = R0_en & R0_addr_sel == 8'h8d;
  assign mem_141_1_W0_addr = W0_addr[25:0];
  assign mem_141_1_W0_clk = W0_clk;
  assign mem_141_1_W0_data = W0_data[15:8];
  assign mem_141_1_W0_en = W0_en & W0_addr_sel == 8'h8d;
  assign mem_141_1_W0_mask = W0_mask[1];
  assign mem_141_2_R0_addr = R0_addr[25:0];
  assign mem_141_2_R0_clk = R0_clk;
  assign mem_141_2_R0_en = R0_en & R0_addr_sel == 8'h8d;
  assign mem_141_2_W0_addr = W0_addr[25:0];
  assign mem_141_2_W0_clk = W0_clk;
  assign mem_141_2_W0_data = W0_data[23:16];
  assign mem_141_2_W0_en = W0_en & W0_addr_sel == 8'h8d;
  assign mem_141_2_W0_mask = W0_mask[2];
  assign mem_141_3_R0_addr = R0_addr[25:0];
  assign mem_141_3_R0_clk = R0_clk;
  assign mem_141_3_R0_en = R0_en & R0_addr_sel == 8'h8d;
  assign mem_141_3_W0_addr = W0_addr[25:0];
  assign mem_141_3_W0_clk = W0_clk;
  assign mem_141_3_W0_data = W0_data[31:24];
  assign mem_141_3_W0_en = W0_en & W0_addr_sel == 8'h8d;
  assign mem_141_3_W0_mask = W0_mask[3];
  assign mem_141_4_R0_addr = R0_addr[25:0];
  assign mem_141_4_R0_clk = R0_clk;
  assign mem_141_4_R0_en = R0_en & R0_addr_sel == 8'h8d;
  assign mem_141_4_W0_addr = W0_addr[25:0];
  assign mem_141_4_W0_clk = W0_clk;
  assign mem_141_4_W0_data = W0_data[39:32];
  assign mem_141_4_W0_en = W0_en & W0_addr_sel == 8'h8d;
  assign mem_141_4_W0_mask = W0_mask[4];
  assign mem_141_5_R0_addr = R0_addr[25:0];
  assign mem_141_5_R0_clk = R0_clk;
  assign mem_141_5_R0_en = R0_en & R0_addr_sel == 8'h8d;
  assign mem_141_5_W0_addr = W0_addr[25:0];
  assign mem_141_5_W0_clk = W0_clk;
  assign mem_141_5_W0_data = W0_data[47:40];
  assign mem_141_5_W0_en = W0_en & W0_addr_sel == 8'h8d;
  assign mem_141_5_W0_mask = W0_mask[5];
  assign mem_141_6_R0_addr = R0_addr[25:0];
  assign mem_141_6_R0_clk = R0_clk;
  assign mem_141_6_R0_en = R0_en & R0_addr_sel == 8'h8d;
  assign mem_141_6_W0_addr = W0_addr[25:0];
  assign mem_141_6_W0_clk = W0_clk;
  assign mem_141_6_W0_data = W0_data[55:48];
  assign mem_141_6_W0_en = W0_en & W0_addr_sel == 8'h8d;
  assign mem_141_6_W0_mask = W0_mask[6];
  assign mem_141_7_R0_addr = R0_addr[25:0];
  assign mem_141_7_R0_clk = R0_clk;
  assign mem_141_7_R0_en = R0_en & R0_addr_sel == 8'h8d;
  assign mem_141_7_W0_addr = W0_addr[25:0];
  assign mem_141_7_W0_clk = W0_clk;
  assign mem_141_7_W0_data = W0_data[63:56];
  assign mem_141_7_W0_en = W0_en & W0_addr_sel == 8'h8d;
  assign mem_141_7_W0_mask = W0_mask[7];
  assign mem_142_0_R0_addr = R0_addr[25:0];
  assign mem_142_0_R0_clk = R0_clk;
  assign mem_142_0_R0_en = R0_en & R0_addr_sel == 8'h8e;
  assign mem_142_0_W0_addr = W0_addr[25:0];
  assign mem_142_0_W0_clk = W0_clk;
  assign mem_142_0_W0_data = W0_data[7:0];
  assign mem_142_0_W0_en = W0_en & W0_addr_sel == 8'h8e;
  assign mem_142_0_W0_mask = W0_mask[0];
  assign mem_142_1_R0_addr = R0_addr[25:0];
  assign mem_142_1_R0_clk = R0_clk;
  assign mem_142_1_R0_en = R0_en & R0_addr_sel == 8'h8e;
  assign mem_142_1_W0_addr = W0_addr[25:0];
  assign mem_142_1_W0_clk = W0_clk;
  assign mem_142_1_W0_data = W0_data[15:8];
  assign mem_142_1_W0_en = W0_en & W0_addr_sel == 8'h8e;
  assign mem_142_1_W0_mask = W0_mask[1];
  assign mem_142_2_R0_addr = R0_addr[25:0];
  assign mem_142_2_R0_clk = R0_clk;
  assign mem_142_2_R0_en = R0_en & R0_addr_sel == 8'h8e;
  assign mem_142_2_W0_addr = W0_addr[25:0];
  assign mem_142_2_W0_clk = W0_clk;
  assign mem_142_2_W0_data = W0_data[23:16];
  assign mem_142_2_W0_en = W0_en & W0_addr_sel == 8'h8e;
  assign mem_142_2_W0_mask = W0_mask[2];
  assign mem_142_3_R0_addr = R0_addr[25:0];
  assign mem_142_3_R0_clk = R0_clk;
  assign mem_142_3_R0_en = R0_en & R0_addr_sel == 8'h8e;
  assign mem_142_3_W0_addr = W0_addr[25:0];
  assign mem_142_3_W0_clk = W0_clk;
  assign mem_142_3_W0_data = W0_data[31:24];
  assign mem_142_3_W0_en = W0_en & W0_addr_sel == 8'h8e;
  assign mem_142_3_W0_mask = W0_mask[3];
  assign mem_142_4_R0_addr = R0_addr[25:0];
  assign mem_142_4_R0_clk = R0_clk;
  assign mem_142_4_R0_en = R0_en & R0_addr_sel == 8'h8e;
  assign mem_142_4_W0_addr = W0_addr[25:0];
  assign mem_142_4_W0_clk = W0_clk;
  assign mem_142_4_W0_data = W0_data[39:32];
  assign mem_142_4_W0_en = W0_en & W0_addr_sel == 8'h8e;
  assign mem_142_4_W0_mask = W0_mask[4];
  assign mem_142_5_R0_addr = R0_addr[25:0];
  assign mem_142_5_R0_clk = R0_clk;
  assign mem_142_5_R0_en = R0_en & R0_addr_sel == 8'h8e;
  assign mem_142_5_W0_addr = W0_addr[25:0];
  assign mem_142_5_W0_clk = W0_clk;
  assign mem_142_5_W0_data = W0_data[47:40];
  assign mem_142_5_W0_en = W0_en & W0_addr_sel == 8'h8e;
  assign mem_142_5_W0_mask = W0_mask[5];
  assign mem_142_6_R0_addr = R0_addr[25:0];
  assign mem_142_6_R0_clk = R0_clk;
  assign mem_142_6_R0_en = R0_en & R0_addr_sel == 8'h8e;
  assign mem_142_6_W0_addr = W0_addr[25:0];
  assign mem_142_6_W0_clk = W0_clk;
  assign mem_142_6_W0_data = W0_data[55:48];
  assign mem_142_6_W0_en = W0_en & W0_addr_sel == 8'h8e;
  assign mem_142_6_W0_mask = W0_mask[6];
  assign mem_142_7_R0_addr = R0_addr[25:0];
  assign mem_142_7_R0_clk = R0_clk;
  assign mem_142_7_R0_en = R0_en & R0_addr_sel == 8'h8e;
  assign mem_142_7_W0_addr = W0_addr[25:0];
  assign mem_142_7_W0_clk = W0_clk;
  assign mem_142_7_W0_data = W0_data[63:56];
  assign mem_142_7_W0_en = W0_en & W0_addr_sel == 8'h8e;
  assign mem_142_7_W0_mask = W0_mask[7];
  assign mem_143_0_R0_addr = R0_addr[25:0];
  assign mem_143_0_R0_clk = R0_clk;
  assign mem_143_0_R0_en = R0_en & R0_addr_sel == 8'h8f;
  assign mem_143_0_W0_addr = W0_addr[25:0];
  assign mem_143_0_W0_clk = W0_clk;
  assign mem_143_0_W0_data = W0_data[7:0];
  assign mem_143_0_W0_en = W0_en & W0_addr_sel == 8'h8f;
  assign mem_143_0_W0_mask = W0_mask[0];
  assign mem_143_1_R0_addr = R0_addr[25:0];
  assign mem_143_1_R0_clk = R0_clk;
  assign mem_143_1_R0_en = R0_en & R0_addr_sel == 8'h8f;
  assign mem_143_1_W0_addr = W0_addr[25:0];
  assign mem_143_1_W0_clk = W0_clk;
  assign mem_143_1_W0_data = W0_data[15:8];
  assign mem_143_1_W0_en = W0_en & W0_addr_sel == 8'h8f;
  assign mem_143_1_W0_mask = W0_mask[1];
  assign mem_143_2_R0_addr = R0_addr[25:0];
  assign mem_143_2_R0_clk = R0_clk;
  assign mem_143_2_R0_en = R0_en & R0_addr_sel == 8'h8f;
  assign mem_143_2_W0_addr = W0_addr[25:0];
  assign mem_143_2_W0_clk = W0_clk;
  assign mem_143_2_W0_data = W0_data[23:16];
  assign mem_143_2_W0_en = W0_en & W0_addr_sel == 8'h8f;
  assign mem_143_2_W0_mask = W0_mask[2];
  assign mem_143_3_R0_addr = R0_addr[25:0];
  assign mem_143_3_R0_clk = R0_clk;
  assign mem_143_3_R0_en = R0_en & R0_addr_sel == 8'h8f;
  assign mem_143_3_W0_addr = W0_addr[25:0];
  assign mem_143_3_W0_clk = W0_clk;
  assign mem_143_3_W0_data = W0_data[31:24];
  assign mem_143_3_W0_en = W0_en & W0_addr_sel == 8'h8f;
  assign mem_143_3_W0_mask = W0_mask[3];
  assign mem_143_4_R0_addr = R0_addr[25:0];
  assign mem_143_4_R0_clk = R0_clk;
  assign mem_143_4_R0_en = R0_en & R0_addr_sel == 8'h8f;
  assign mem_143_4_W0_addr = W0_addr[25:0];
  assign mem_143_4_W0_clk = W0_clk;
  assign mem_143_4_W0_data = W0_data[39:32];
  assign mem_143_4_W0_en = W0_en & W0_addr_sel == 8'h8f;
  assign mem_143_4_W0_mask = W0_mask[4];
  assign mem_143_5_R0_addr = R0_addr[25:0];
  assign mem_143_5_R0_clk = R0_clk;
  assign mem_143_5_R0_en = R0_en & R0_addr_sel == 8'h8f;
  assign mem_143_5_W0_addr = W0_addr[25:0];
  assign mem_143_5_W0_clk = W0_clk;
  assign mem_143_5_W0_data = W0_data[47:40];
  assign mem_143_5_W0_en = W0_en & W0_addr_sel == 8'h8f;
  assign mem_143_5_W0_mask = W0_mask[5];
  assign mem_143_6_R0_addr = R0_addr[25:0];
  assign mem_143_6_R0_clk = R0_clk;
  assign mem_143_6_R0_en = R0_en & R0_addr_sel == 8'h8f;
  assign mem_143_6_W0_addr = W0_addr[25:0];
  assign mem_143_6_W0_clk = W0_clk;
  assign mem_143_6_W0_data = W0_data[55:48];
  assign mem_143_6_W0_en = W0_en & W0_addr_sel == 8'h8f;
  assign mem_143_6_W0_mask = W0_mask[6];
  assign mem_143_7_R0_addr = R0_addr[25:0];
  assign mem_143_7_R0_clk = R0_clk;
  assign mem_143_7_R0_en = R0_en & R0_addr_sel == 8'h8f;
  assign mem_143_7_W0_addr = W0_addr[25:0];
  assign mem_143_7_W0_clk = W0_clk;
  assign mem_143_7_W0_data = W0_data[63:56];
  assign mem_143_7_W0_en = W0_en & W0_addr_sel == 8'h8f;
  assign mem_143_7_W0_mask = W0_mask[7];
  assign mem_144_0_R0_addr = R0_addr[25:0];
  assign mem_144_0_R0_clk = R0_clk;
  assign mem_144_0_R0_en = R0_en & R0_addr_sel == 8'h90;
  assign mem_144_0_W0_addr = W0_addr[25:0];
  assign mem_144_0_W0_clk = W0_clk;
  assign mem_144_0_W0_data = W0_data[7:0];
  assign mem_144_0_W0_en = W0_en & W0_addr_sel == 8'h90;
  assign mem_144_0_W0_mask = W0_mask[0];
  assign mem_144_1_R0_addr = R0_addr[25:0];
  assign mem_144_1_R0_clk = R0_clk;
  assign mem_144_1_R0_en = R0_en & R0_addr_sel == 8'h90;
  assign mem_144_1_W0_addr = W0_addr[25:0];
  assign mem_144_1_W0_clk = W0_clk;
  assign mem_144_1_W0_data = W0_data[15:8];
  assign mem_144_1_W0_en = W0_en & W0_addr_sel == 8'h90;
  assign mem_144_1_W0_mask = W0_mask[1];
  assign mem_144_2_R0_addr = R0_addr[25:0];
  assign mem_144_2_R0_clk = R0_clk;
  assign mem_144_2_R0_en = R0_en & R0_addr_sel == 8'h90;
  assign mem_144_2_W0_addr = W0_addr[25:0];
  assign mem_144_2_W0_clk = W0_clk;
  assign mem_144_2_W0_data = W0_data[23:16];
  assign mem_144_2_W0_en = W0_en & W0_addr_sel == 8'h90;
  assign mem_144_2_W0_mask = W0_mask[2];
  assign mem_144_3_R0_addr = R0_addr[25:0];
  assign mem_144_3_R0_clk = R0_clk;
  assign mem_144_3_R0_en = R0_en & R0_addr_sel == 8'h90;
  assign mem_144_3_W0_addr = W0_addr[25:0];
  assign mem_144_3_W0_clk = W0_clk;
  assign mem_144_3_W0_data = W0_data[31:24];
  assign mem_144_3_W0_en = W0_en & W0_addr_sel == 8'h90;
  assign mem_144_3_W0_mask = W0_mask[3];
  assign mem_144_4_R0_addr = R0_addr[25:0];
  assign mem_144_4_R0_clk = R0_clk;
  assign mem_144_4_R0_en = R0_en & R0_addr_sel == 8'h90;
  assign mem_144_4_W0_addr = W0_addr[25:0];
  assign mem_144_4_W0_clk = W0_clk;
  assign mem_144_4_W0_data = W0_data[39:32];
  assign mem_144_4_W0_en = W0_en & W0_addr_sel == 8'h90;
  assign mem_144_4_W0_mask = W0_mask[4];
  assign mem_144_5_R0_addr = R0_addr[25:0];
  assign mem_144_5_R0_clk = R0_clk;
  assign mem_144_5_R0_en = R0_en & R0_addr_sel == 8'h90;
  assign mem_144_5_W0_addr = W0_addr[25:0];
  assign mem_144_5_W0_clk = W0_clk;
  assign mem_144_5_W0_data = W0_data[47:40];
  assign mem_144_5_W0_en = W0_en & W0_addr_sel == 8'h90;
  assign mem_144_5_W0_mask = W0_mask[5];
  assign mem_144_6_R0_addr = R0_addr[25:0];
  assign mem_144_6_R0_clk = R0_clk;
  assign mem_144_6_R0_en = R0_en & R0_addr_sel == 8'h90;
  assign mem_144_6_W0_addr = W0_addr[25:0];
  assign mem_144_6_W0_clk = W0_clk;
  assign mem_144_6_W0_data = W0_data[55:48];
  assign mem_144_6_W0_en = W0_en & W0_addr_sel == 8'h90;
  assign mem_144_6_W0_mask = W0_mask[6];
  assign mem_144_7_R0_addr = R0_addr[25:0];
  assign mem_144_7_R0_clk = R0_clk;
  assign mem_144_7_R0_en = R0_en & R0_addr_sel == 8'h90;
  assign mem_144_7_W0_addr = W0_addr[25:0];
  assign mem_144_7_W0_clk = W0_clk;
  assign mem_144_7_W0_data = W0_data[63:56];
  assign mem_144_7_W0_en = W0_en & W0_addr_sel == 8'h90;
  assign mem_144_7_W0_mask = W0_mask[7];
  assign mem_145_0_R0_addr = R0_addr[25:0];
  assign mem_145_0_R0_clk = R0_clk;
  assign mem_145_0_R0_en = R0_en & R0_addr_sel == 8'h91;
  assign mem_145_0_W0_addr = W0_addr[25:0];
  assign mem_145_0_W0_clk = W0_clk;
  assign mem_145_0_W0_data = W0_data[7:0];
  assign mem_145_0_W0_en = W0_en & W0_addr_sel == 8'h91;
  assign mem_145_0_W0_mask = W0_mask[0];
  assign mem_145_1_R0_addr = R0_addr[25:0];
  assign mem_145_1_R0_clk = R0_clk;
  assign mem_145_1_R0_en = R0_en & R0_addr_sel == 8'h91;
  assign mem_145_1_W0_addr = W0_addr[25:0];
  assign mem_145_1_W0_clk = W0_clk;
  assign mem_145_1_W0_data = W0_data[15:8];
  assign mem_145_1_W0_en = W0_en & W0_addr_sel == 8'h91;
  assign mem_145_1_W0_mask = W0_mask[1];
  assign mem_145_2_R0_addr = R0_addr[25:0];
  assign mem_145_2_R0_clk = R0_clk;
  assign mem_145_2_R0_en = R0_en & R0_addr_sel == 8'h91;
  assign mem_145_2_W0_addr = W0_addr[25:0];
  assign mem_145_2_W0_clk = W0_clk;
  assign mem_145_2_W0_data = W0_data[23:16];
  assign mem_145_2_W0_en = W0_en & W0_addr_sel == 8'h91;
  assign mem_145_2_W0_mask = W0_mask[2];
  assign mem_145_3_R0_addr = R0_addr[25:0];
  assign mem_145_3_R0_clk = R0_clk;
  assign mem_145_3_R0_en = R0_en & R0_addr_sel == 8'h91;
  assign mem_145_3_W0_addr = W0_addr[25:0];
  assign mem_145_3_W0_clk = W0_clk;
  assign mem_145_3_W0_data = W0_data[31:24];
  assign mem_145_3_W0_en = W0_en & W0_addr_sel == 8'h91;
  assign mem_145_3_W0_mask = W0_mask[3];
  assign mem_145_4_R0_addr = R0_addr[25:0];
  assign mem_145_4_R0_clk = R0_clk;
  assign mem_145_4_R0_en = R0_en & R0_addr_sel == 8'h91;
  assign mem_145_4_W0_addr = W0_addr[25:0];
  assign mem_145_4_W0_clk = W0_clk;
  assign mem_145_4_W0_data = W0_data[39:32];
  assign mem_145_4_W0_en = W0_en & W0_addr_sel == 8'h91;
  assign mem_145_4_W0_mask = W0_mask[4];
  assign mem_145_5_R0_addr = R0_addr[25:0];
  assign mem_145_5_R0_clk = R0_clk;
  assign mem_145_5_R0_en = R0_en & R0_addr_sel == 8'h91;
  assign mem_145_5_W0_addr = W0_addr[25:0];
  assign mem_145_5_W0_clk = W0_clk;
  assign mem_145_5_W0_data = W0_data[47:40];
  assign mem_145_5_W0_en = W0_en & W0_addr_sel == 8'h91;
  assign mem_145_5_W0_mask = W0_mask[5];
  assign mem_145_6_R0_addr = R0_addr[25:0];
  assign mem_145_6_R0_clk = R0_clk;
  assign mem_145_6_R0_en = R0_en & R0_addr_sel == 8'h91;
  assign mem_145_6_W0_addr = W0_addr[25:0];
  assign mem_145_6_W0_clk = W0_clk;
  assign mem_145_6_W0_data = W0_data[55:48];
  assign mem_145_6_W0_en = W0_en & W0_addr_sel == 8'h91;
  assign mem_145_6_W0_mask = W0_mask[6];
  assign mem_145_7_R0_addr = R0_addr[25:0];
  assign mem_145_7_R0_clk = R0_clk;
  assign mem_145_7_R0_en = R0_en & R0_addr_sel == 8'h91;
  assign mem_145_7_W0_addr = W0_addr[25:0];
  assign mem_145_7_W0_clk = W0_clk;
  assign mem_145_7_W0_data = W0_data[63:56];
  assign mem_145_7_W0_en = W0_en & W0_addr_sel == 8'h91;
  assign mem_145_7_W0_mask = W0_mask[7];
  assign mem_146_0_R0_addr = R0_addr[25:0];
  assign mem_146_0_R0_clk = R0_clk;
  assign mem_146_0_R0_en = R0_en & R0_addr_sel == 8'h92;
  assign mem_146_0_W0_addr = W0_addr[25:0];
  assign mem_146_0_W0_clk = W0_clk;
  assign mem_146_0_W0_data = W0_data[7:0];
  assign mem_146_0_W0_en = W0_en & W0_addr_sel == 8'h92;
  assign mem_146_0_W0_mask = W0_mask[0];
  assign mem_146_1_R0_addr = R0_addr[25:0];
  assign mem_146_1_R0_clk = R0_clk;
  assign mem_146_1_R0_en = R0_en & R0_addr_sel == 8'h92;
  assign mem_146_1_W0_addr = W0_addr[25:0];
  assign mem_146_1_W0_clk = W0_clk;
  assign mem_146_1_W0_data = W0_data[15:8];
  assign mem_146_1_W0_en = W0_en & W0_addr_sel == 8'h92;
  assign mem_146_1_W0_mask = W0_mask[1];
  assign mem_146_2_R0_addr = R0_addr[25:0];
  assign mem_146_2_R0_clk = R0_clk;
  assign mem_146_2_R0_en = R0_en & R0_addr_sel == 8'h92;
  assign mem_146_2_W0_addr = W0_addr[25:0];
  assign mem_146_2_W0_clk = W0_clk;
  assign mem_146_2_W0_data = W0_data[23:16];
  assign mem_146_2_W0_en = W0_en & W0_addr_sel == 8'h92;
  assign mem_146_2_W0_mask = W0_mask[2];
  assign mem_146_3_R0_addr = R0_addr[25:0];
  assign mem_146_3_R0_clk = R0_clk;
  assign mem_146_3_R0_en = R0_en & R0_addr_sel == 8'h92;
  assign mem_146_3_W0_addr = W0_addr[25:0];
  assign mem_146_3_W0_clk = W0_clk;
  assign mem_146_3_W0_data = W0_data[31:24];
  assign mem_146_3_W0_en = W0_en & W0_addr_sel == 8'h92;
  assign mem_146_3_W0_mask = W0_mask[3];
  assign mem_146_4_R0_addr = R0_addr[25:0];
  assign mem_146_4_R0_clk = R0_clk;
  assign mem_146_4_R0_en = R0_en & R0_addr_sel == 8'h92;
  assign mem_146_4_W0_addr = W0_addr[25:0];
  assign mem_146_4_W0_clk = W0_clk;
  assign mem_146_4_W0_data = W0_data[39:32];
  assign mem_146_4_W0_en = W0_en & W0_addr_sel == 8'h92;
  assign mem_146_4_W0_mask = W0_mask[4];
  assign mem_146_5_R0_addr = R0_addr[25:0];
  assign mem_146_5_R0_clk = R0_clk;
  assign mem_146_5_R0_en = R0_en & R0_addr_sel == 8'h92;
  assign mem_146_5_W0_addr = W0_addr[25:0];
  assign mem_146_5_W0_clk = W0_clk;
  assign mem_146_5_W0_data = W0_data[47:40];
  assign mem_146_5_W0_en = W0_en & W0_addr_sel == 8'h92;
  assign mem_146_5_W0_mask = W0_mask[5];
  assign mem_146_6_R0_addr = R0_addr[25:0];
  assign mem_146_6_R0_clk = R0_clk;
  assign mem_146_6_R0_en = R0_en & R0_addr_sel == 8'h92;
  assign mem_146_6_W0_addr = W0_addr[25:0];
  assign mem_146_6_W0_clk = W0_clk;
  assign mem_146_6_W0_data = W0_data[55:48];
  assign mem_146_6_W0_en = W0_en & W0_addr_sel == 8'h92;
  assign mem_146_6_W0_mask = W0_mask[6];
  assign mem_146_7_R0_addr = R0_addr[25:0];
  assign mem_146_7_R0_clk = R0_clk;
  assign mem_146_7_R0_en = R0_en & R0_addr_sel == 8'h92;
  assign mem_146_7_W0_addr = W0_addr[25:0];
  assign mem_146_7_W0_clk = W0_clk;
  assign mem_146_7_W0_data = W0_data[63:56];
  assign mem_146_7_W0_en = W0_en & W0_addr_sel == 8'h92;
  assign mem_146_7_W0_mask = W0_mask[7];
  assign mem_147_0_R0_addr = R0_addr[25:0];
  assign mem_147_0_R0_clk = R0_clk;
  assign mem_147_0_R0_en = R0_en & R0_addr_sel == 8'h93;
  assign mem_147_0_W0_addr = W0_addr[25:0];
  assign mem_147_0_W0_clk = W0_clk;
  assign mem_147_0_W0_data = W0_data[7:0];
  assign mem_147_0_W0_en = W0_en & W0_addr_sel == 8'h93;
  assign mem_147_0_W0_mask = W0_mask[0];
  assign mem_147_1_R0_addr = R0_addr[25:0];
  assign mem_147_1_R0_clk = R0_clk;
  assign mem_147_1_R0_en = R0_en & R0_addr_sel == 8'h93;
  assign mem_147_1_W0_addr = W0_addr[25:0];
  assign mem_147_1_W0_clk = W0_clk;
  assign mem_147_1_W0_data = W0_data[15:8];
  assign mem_147_1_W0_en = W0_en & W0_addr_sel == 8'h93;
  assign mem_147_1_W0_mask = W0_mask[1];
  assign mem_147_2_R0_addr = R0_addr[25:0];
  assign mem_147_2_R0_clk = R0_clk;
  assign mem_147_2_R0_en = R0_en & R0_addr_sel == 8'h93;
  assign mem_147_2_W0_addr = W0_addr[25:0];
  assign mem_147_2_W0_clk = W0_clk;
  assign mem_147_2_W0_data = W0_data[23:16];
  assign mem_147_2_W0_en = W0_en & W0_addr_sel == 8'h93;
  assign mem_147_2_W0_mask = W0_mask[2];
  assign mem_147_3_R0_addr = R0_addr[25:0];
  assign mem_147_3_R0_clk = R0_clk;
  assign mem_147_3_R0_en = R0_en & R0_addr_sel == 8'h93;
  assign mem_147_3_W0_addr = W0_addr[25:0];
  assign mem_147_3_W0_clk = W0_clk;
  assign mem_147_3_W0_data = W0_data[31:24];
  assign mem_147_3_W0_en = W0_en & W0_addr_sel == 8'h93;
  assign mem_147_3_W0_mask = W0_mask[3];
  assign mem_147_4_R0_addr = R0_addr[25:0];
  assign mem_147_4_R0_clk = R0_clk;
  assign mem_147_4_R0_en = R0_en & R0_addr_sel == 8'h93;
  assign mem_147_4_W0_addr = W0_addr[25:0];
  assign mem_147_4_W0_clk = W0_clk;
  assign mem_147_4_W0_data = W0_data[39:32];
  assign mem_147_4_W0_en = W0_en & W0_addr_sel == 8'h93;
  assign mem_147_4_W0_mask = W0_mask[4];
  assign mem_147_5_R0_addr = R0_addr[25:0];
  assign mem_147_5_R0_clk = R0_clk;
  assign mem_147_5_R0_en = R0_en & R0_addr_sel == 8'h93;
  assign mem_147_5_W0_addr = W0_addr[25:0];
  assign mem_147_5_W0_clk = W0_clk;
  assign mem_147_5_W0_data = W0_data[47:40];
  assign mem_147_5_W0_en = W0_en & W0_addr_sel == 8'h93;
  assign mem_147_5_W0_mask = W0_mask[5];
  assign mem_147_6_R0_addr = R0_addr[25:0];
  assign mem_147_6_R0_clk = R0_clk;
  assign mem_147_6_R0_en = R0_en & R0_addr_sel == 8'h93;
  assign mem_147_6_W0_addr = W0_addr[25:0];
  assign mem_147_6_W0_clk = W0_clk;
  assign mem_147_6_W0_data = W0_data[55:48];
  assign mem_147_6_W0_en = W0_en & W0_addr_sel == 8'h93;
  assign mem_147_6_W0_mask = W0_mask[6];
  assign mem_147_7_R0_addr = R0_addr[25:0];
  assign mem_147_7_R0_clk = R0_clk;
  assign mem_147_7_R0_en = R0_en & R0_addr_sel == 8'h93;
  assign mem_147_7_W0_addr = W0_addr[25:0];
  assign mem_147_7_W0_clk = W0_clk;
  assign mem_147_7_W0_data = W0_data[63:56];
  assign mem_147_7_W0_en = W0_en & W0_addr_sel == 8'h93;
  assign mem_147_7_W0_mask = W0_mask[7];
  assign mem_148_0_R0_addr = R0_addr[25:0];
  assign mem_148_0_R0_clk = R0_clk;
  assign mem_148_0_R0_en = R0_en & R0_addr_sel == 8'h94;
  assign mem_148_0_W0_addr = W0_addr[25:0];
  assign mem_148_0_W0_clk = W0_clk;
  assign mem_148_0_W0_data = W0_data[7:0];
  assign mem_148_0_W0_en = W0_en & W0_addr_sel == 8'h94;
  assign mem_148_0_W0_mask = W0_mask[0];
  assign mem_148_1_R0_addr = R0_addr[25:0];
  assign mem_148_1_R0_clk = R0_clk;
  assign mem_148_1_R0_en = R0_en & R0_addr_sel == 8'h94;
  assign mem_148_1_W0_addr = W0_addr[25:0];
  assign mem_148_1_W0_clk = W0_clk;
  assign mem_148_1_W0_data = W0_data[15:8];
  assign mem_148_1_W0_en = W0_en & W0_addr_sel == 8'h94;
  assign mem_148_1_W0_mask = W0_mask[1];
  assign mem_148_2_R0_addr = R0_addr[25:0];
  assign mem_148_2_R0_clk = R0_clk;
  assign mem_148_2_R0_en = R0_en & R0_addr_sel == 8'h94;
  assign mem_148_2_W0_addr = W0_addr[25:0];
  assign mem_148_2_W0_clk = W0_clk;
  assign mem_148_2_W0_data = W0_data[23:16];
  assign mem_148_2_W0_en = W0_en & W0_addr_sel == 8'h94;
  assign mem_148_2_W0_mask = W0_mask[2];
  assign mem_148_3_R0_addr = R0_addr[25:0];
  assign mem_148_3_R0_clk = R0_clk;
  assign mem_148_3_R0_en = R0_en & R0_addr_sel == 8'h94;
  assign mem_148_3_W0_addr = W0_addr[25:0];
  assign mem_148_3_W0_clk = W0_clk;
  assign mem_148_3_W0_data = W0_data[31:24];
  assign mem_148_3_W0_en = W0_en & W0_addr_sel == 8'h94;
  assign mem_148_3_W0_mask = W0_mask[3];
  assign mem_148_4_R0_addr = R0_addr[25:0];
  assign mem_148_4_R0_clk = R0_clk;
  assign mem_148_4_R0_en = R0_en & R0_addr_sel == 8'h94;
  assign mem_148_4_W0_addr = W0_addr[25:0];
  assign mem_148_4_W0_clk = W0_clk;
  assign mem_148_4_W0_data = W0_data[39:32];
  assign mem_148_4_W0_en = W0_en & W0_addr_sel == 8'h94;
  assign mem_148_4_W0_mask = W0_mask[4];
  assign mem_148_5_R0_addr = R0_addr[25:0];
  assign mem_148_5_R0_clk = R0_clk;
  assign mem_148_5_R0_en = R0_en & R0_addr_sel == 8'h94;
  assign mem_148_5_W0_addr = W0_addr[25:0];
  assign mem_148_5_W0_clk = W0_clk;
  assign mem_148_5_W0_data = W0_data[47:40];
  assign mem_148_5_W0_en = W0_en & W0_addr_sel == 8'h94;
  assign mem_148_5_W0_mask = W0_mask[5];
  assign mem_148_6_R0_addr = R0_addr[25:0];
  assign mem_148_6_R0_clk = R0_clk;
  assign mem_148_6_R0_en = R0_en & R0_addr_sel == 8'h94;
  assign mem_148_6_W0_addr = W0_addr[25:0];
  assign mem_148_6_W0_clk = W0_clk;
  assign mem_148_6_W0_data = W0_data[55:48];
  assign mem_148_6_W0_en = W0_en & W0_addr_sel == 8'h94;
  assign mem_148_6_W0_mask = W0_mask[6];
  assign mem_148_7_R0_addr = R0_addr[25:0];
  assign mem_148_7_R0_clk = R0_clk;
  assign mem_148_7_R0_en = R0_en & R0_addr_sel == 8'h94;
  assign mem_148_7_W0_addr = W0_addr[25:0];
  assign mem_148_7_W0_clk = W0_clk;
  assign mem_148_7_W0_data = W0_data[63:56];
  assign mem_148_7_W0_en = W0_en & W0_addr_sel == 8'h94;
  assign mem_148_7_W0_mask = W0_mask[7];
  assign mem_149_0_R0_addr = R0_addr[25:0];
  assign mem_149_0_R0_clk = R0_clk;
  assign mem_149_0_R0_en = R0_en & R0_addr_sel == 8'h95;
  assign mem_149_0_W0_addr = W0_addr[25:0];
  assign mem_149_0_W0_clk = W0_clk;
  assign mem_149_0_W0_data = W0_data[7:0];
  assign mem_149_0_W0_en = W0_en & W0_addr_sel == 8'h95;
  assign mem_149_0_W0_mask = W0_mask[0];
  assign mem_149_1_R0_addr = R0_addr[25:0];
  assign mem_149_1_R0_clk = R0_clk;
  assign mem_149_1_R0_en = R0_en & R0_addr_sel == 8'h95;
  assign mem_149_1_W0_addr = W0_addr[25:0];
  assign mem_149_1_W0_clk = W0_clk;
  assign mem_149_1_W0_data = W0_data[15:8];
  assign mem_149_1_W0_en = W0_en & W0_addr_sel == 8'h95;
  assign mem_149_1_W0_mask = W0_mask[1];
  assign mem_149_2_R0_addr = R0_addr[25:0];
  assign mem_149_2_R0_clk = R0_clk;
  assign mem_149_2_R0_en = R0_en & R0_addr_sel == 8'h95;
  assign mem_149_2_W0_addr = W0_addr[25:0];
  assign mem_149_2_W0_clk = W0_clk;
  assign mem_149_2_W0_data = W0_data[23:16];
  assign mem_149_2_W0_en = W0_en & W0_addr_sel == 8'h95;
  assign mem_149_2_W0_mask = W0_mask[2];
  assign mem_149_3_R0_addr = R0_addr[25:0];
  assign mem_149_3_R0_clk = R0_clk;
  assign mem_149_3_R0_en = R0_en & R0_addr_sel == 8'h95;
  assign mem_149_3_W0_addr = W0_addr[25:0];
  assign mem_149_3_W0_clk = W0_clk;
  assign mem_149_3_W0_data = W0_data[31:24];
  assign mem_149_3_W0_en = W0_en & W0_addr_sel == 8'h95;
  assign mem_149_3_W0_mask = W0_mask[3];
  assign mem_149_4_R0_addr = R0_addr[25:0];
  assign mem_149_4_R0_clk = R0_clk;
  assign mem_149_4_R0_en = R0_en & R0_addr_sel == 8'h95;
  assign mem_149_4_W0_addr = W0_addr[25:0];
  assign mem_149_4_W0_clk = W0_clk;
  assign mem_149_4_W0_data = W0_data[39:32];
  assign mem_149_4_W0_en = W0_en & W0_addr_sel == 8'h95;
  assign mem_149_4_W0_mask = W0_mask[4];
  assign mem_149_5_R0_addr = R0_addr[25:0];
  assign mem_149_5_R0_clk = R0_clk;
  assign mem_149_5_R0_en = R0_en & R0_addr_sel == 8'h95;
  assign mem_149_5_W0_addr = W0_addr[25:0];
  assign mem_149_5_W0_clk = W0_clk;
  assign mem_149_5_W0_data = W0_data[47:40];
  assign mem_149_5_W0_en = W0_en & W0_addr_sel == 8'h95;
  assign mem_149_5_W0_mask = W0_mask[5];
  assign mem_149_6_R0_addr = R0_addr[25:0];
  assign mem_149_6_R0_clk = R0_clk;
  assign mem_149_6_R0_en = R0_en & R0_addr_sel == 8'h95;
  assign mem_149_6_W0_addr = W0_addr[25:0];
  assign mem_149_6_W0_clk = W0_clk;
  assign mem_149_6_W0_data = W0_data[55:48];
  assign mem_149_6_W0_en = W0_en & W0_addr_sel == 8'h95;
  assign mem_149_6_W0_mask = W0_mask[6];
  assign mem_149_7_R0_addr = R0_addr[25:0];
  assign mem_149_7_R0_clk = R0_clk;
  assign mem_149_7_R0_en = R0_en & R0_addr_sel == 8'h95;
  assign mem_149_7_W0_addr = W0_addr[25:0];
  assign mem_149_7_W0_clk = W0_clk;
  assign mem_149_7_W0_data = W0_data[63:56];
  assign mem_149_7_W0_en = W0_en & W0_addr_sel == 8'h95;
  assign mem_149_7_W0_mask = W0_mask[7];
  assign mem_150_0_R0_addr = R0_addr[25:0];
  assign mem_150_0_R0_clk = R0_clk;
  assign mem_150_0_R0_en = R0_en & R0_addr_sel == 8'h96;
  assign mem_150_0_W0_addr = W0_addr[25:0];
  assign mem_150_0_W0_clk = W0_clk;
  assign mem_150_0_W0_data = W0_data[7:0];
  assign mem_150_0_W0_en = W0_en & W0_addr_sel == 8'h96;
  assign mem_150_0_W0_mask = W0_mask[0];
  assign mem_150_1_R0_addr = R0_addr[25:0];
  assign mem_150_1_R0_clk = R0_clk;
  assign mem_150_1_R0_en = R0_en & R0_addr_sel == 8'h96;
  assign mem_150_1_W0_addr = W0_addr[25:0];
  assign mem_150_1_W0_clk = W0_clk;
  assign mem_150_1_W0_data = W0_data[15:8];
  assign mem_150_1_W0_en = W0_en & W0_addr_sel == 8'h96;
  assign mem_150_1_W0_mask = W0_mask[1];
  assign mem_150_2_R0_addr = R0_addr[25:0];
  assign mem_150_2_R0_clk = R0_clk;
  assign mem_150_2_R0_en = R0_en & R0_addr_sel == 8'h96;
  assign mem_150_2_W0_addr = W0_addr[25:0];
  assign mem_150_2_W0_clk = W0_clk;
  assign mem_150_2_W0_data = W0_data[23:16];
  assign mem_150_2_W0_en = W0_en & W0_addr_sel == 8'h96;
  assign mem_150_2_W0_mask = W0_mask[2];
  assign mem_150_3_R0_addr = R0_addr[25:0];
  assign mem_150_3_R0_clk = R0_clk;
  assign mem_150_3_R0_en = R0_en & R0_addr_sel == 8'h96;
  assign mem_150_3_W0_addr = W0_addr[25:0];
  assign mem_150_3_W0_clk = W0_clk;
  assign mem_150_3_W0_data = W0_data[31:24];
  assign mem_150_3_W0_en = W0_en & W0_addr_sel == 8'h96;
  assign mem_150_3_W0_mask = W0_mask[3];
  assign mem_150_4_R0_addr = R0_addr[25:0];
  assign mem_150_4_R0_clk = R0_clk;
  assign mem_150_4_R0_en = R0_en & R0_addr_sel == 8'h96;
  assign mem_150_4_W0_addr = W0_addr[25:0];
  assign mem_150_4_W0_clk = W0_clk;
  assign mem_150_4_W0_data = W0_data[39:32];
  assign mem_150_4_W0_en = W0_en & W0_addr_sel == 8'h96;
  assign mem_150_4_W0_mask = W0_mask[4];
  assign mem_150_5_R0_addr = R0_addr[25:0];
  assign mem_150_5_R0_clk = R0_clk;
  assign mem_150_5_R0_en = R0_en & R0_addr_sel == 8'h96;
  assign mem_150_5_W0_addr = W0_addr[25:0];
  assign mem_150_5_W0_clk = W0_clk;
  assign mem_150_5_W0_data = W0_data[47:40];
  assign mem_150_5_W0_en = W0_en & W0_addr_sel == 8'h96;
  assign mem_150_5_W0_mask = W0_mask[5];
  assign mem_150_6_R0_addr = R0_addr[25:0];
  assign mem_150_6_R0_clk = R0_clk;
  assign mem_150_6_R0_en = R0_en & R0_addr_sel == 8'h96;
  assign mem_150_6_W0_addr = W0_addr[25:0];
  assign mem_150_6_W0_clk = W0_clk;
  assign mem_150_6_W0_data = W0_data[55:48];
  assign mem_150_6_W0_en = W0_en & W0_addr_sel == 8'h96;
  assign mem_150_6_W0_mask = W0_mask[6];
  assign mem_150_7_R0_addr = R0_addr[25:0];
  assign mem_150_7_R0_clk = R0_clk;
  assign mem_150_7_R0_en = R0_en & R0_addr_sel == 8'h96;
  assign mem_150_7_W0_addr = W0_addr[25:0];
  assign mem_150_7_W0_clk = W0_clk;
  assign mem_150_7_W0_data = W0_data[63:56];
  assign mem_150_7_W0_en = W0_en & W0_addr_sel == 8'h96;
  assign mem_150_7_W0_mask = W0_mask[7];
  assign mem_151_0_R0_addr = R0_addr[25:0];
  assign mem_151_0_R0_clk = R0_clk;
  assign mem_151_0_R0_en = R0_en & R0_addr_sel == 8'h97;
  assign mem_151_0_W0_addr = W0_addr[25:0];
  assign mem_151_0_W0_clk = W0_clk;
  assign mem_151_0_W0_data = W0_data[7:0];
  assign mem_151_0_W0_en = W0_en & W0_addr_sel == 8'h97;
  assign mem_151_0_W0_mask = W0_mask[0];
  assign mem_151_1_R0_addr = R0_addr[25:0];
  assign mem_151_1_R0_clk = R0_clk;
  assign mem_151_1_R0_en = R0_en & R0_addr_sel == 8'h97;
  assign mem_151_1_W0_addr = W0_addr[25:0];
  assign mem_151_1_W0_clk = W0_clk;
  assign mem_151_1_W0_data = W0_data[15:8];
  assign mem_151_1_W0_en = W0_en & W0_addr_sel == 8'h97;
  assign mem_151_1_W0_mask = W0_mask[1];
  assign mem_151_2_R0_addr = R0_addr[25:0];
  assign mem_151_2_R0_clk = R0_clk;
  assign mem_151_2_R0_en = R0_en & R0_addr_sel == 8'h97;
  assign mem_151_2_W0_addr = W0_addr[25:0];
  assign mem_151_2_W0_clk = W0_clk;
  assign mem_151_2_W0_data = W0_data[23:16];
  assign mem_151_2_W0_en = W0_en & W0_addr_sel == 8'h97;
  assign mem_151_2_W0_mask = W0_mask[2];
  assign mem_151_3_R0_addr = R0_addr[25:0];
  assign mem_151_3_R0_clk = R0_clk;
  assign mem_151_3_R0_en = R0_en & R0_addr_sel == 8'h97;
  assign mem_151_3_W0_addr = W0_addr[25:0];
  assign mem_151_3_W0_clk = W0_clk;
  assign mem_151_3_W0_data = W0_data[31:24];
  assign mem_151_3_W0_en = W0_en & W0_addr_sel == 8'h97;
  assign mem_151_3_W0_mask = W0_mask[3];
  assign mem_151_4_R0_addr = R0_addr[25:0];
  assign mem_151_4_R0_clk = R0_clk;
  assign mem_151_4_R0_en = R0_en & R0_addr_sel == 8'h97;
  assign mem_151_4_W0_addr = W0_addr[25:0];
  assign mem_151_4_W0_clk = W0_clk;
  assign mem_151_4_W0_data = W0_data[39:32];
  assign mem_151_4_W0_en = W0_en & W0_addr_sel == 8'h97;
  assign mem_151_4_W0_mask = W0_mask[4];
  assign mem_151_5_R0_addr = R0_addr[25:0];
  assign mem_151_5_R0_clk = R0_clk;
  assign mem_151_5_R0_en = R0_en & R0_addr_sel == 8'h97;
  assign mem_151_5_W0_addr = W0_addr[25:0];
  assign mem_151_5_W0_clk = W0_clk;
  assign mem_151_5_W0_data = W0_data[47:40];
  assign mem_151_5_W0_en = W0_en & W0_addr_sel == 8'h97;
  assign mem_151_5_W0_mask = W0_mask[5];
  assign mem_151_6_R0_addr = R0_addr[25:0];
  assign mem_151_6_R0_clk = R0_clk;
  assign mem_151_6_R0_en = R0_en & R0_addr_sel == 8'h97;
  assign mem_151_6_W0_addr = W0_addr[25:0];
  assign mem_151_6_W0_clk = W0_clk;
  assign mem_151_6_W0_data = W0_data[55:48];
  assign mem_151_6_W0_en = W0_en & W0_addr_sel == 8'h97;
  assign mem_151_6_W0_mask = W0_mask[6];
  assign mem_151_7_R0_addr = R0_addr[25:0];
  assign mem_151_7_R0_clk = R0_clk;
  assign mem_151_7_R0_en = R0_en & R0_addr_sel == 8'h97;
  assign mem_151_7_W0_addr = W0_addr[25:0];
  assign mem_151_7_W0_clk = W0_clk;
  assign mem_151_7_W0_data = W0_data[63:56];
  assign mem_151_7_W0_en = W0_en & W0_addr_sel == 8'h97;
  assign mem_151_7_W0_mask = W0_mask[7];
  assign mem_152_0_R0_addr = R0_addr[25:0];
  assign mem_152_0_R0_clk = R0_clk;
  assign mem_152_0_R0_en = R0_en & R0_addr_sel == 8'h98;
  assign mem_152_0_W0_addr = W0_addr[25:0];
  assign mem_152_0_W0_clk = W0_clk;
  assign mem_152_0_W0_data = W0_data[7:0];
  assign mem_152_0_W0_en = W0_en & W0_addr_sel == 8'h98;
  assign mem_152_0_W0_mask = W0_mask[0];
  assign mem_152_1_R0_addr = R0_addr[25:0];
  assign mem_152_1_R0_clk = R0_clk;
  assign mem_152_1_R0_en = R0_en & R0_addr_sel == 8'h98;
  assign mem_152_1_W0_addr = W0_addr[25:0];
  assign mem_152_1_W0_clk = W0_clk;
  assign mem_152_1_W0_data = W0_data[15:8];
  assign mem_152_1_W0_en = W0_en & W0_addr_sel == 8'h98;
  assign mem_152_1_W0_mask = W0_mask[1];
  assign mem_152_2_R0_addr = R0_addr[25:0];
  assign mem_152_2_R0_clk = R0_clk;
  assign mem_152_2_R0_en = R0_en & R0_addr_sel == 8'h98;
  assign mem_152_2_W0_addr = W0_addr[25:0];
  assign mem_152_2_W0_clk = W0_clk;
  assign mem_152_2_W0_data = W0_data[23:16];
  assign mem_152_2_W0_en = W0_en & W0_addr_sel == 8'h98;
  assign mem_152_2_W0_mask = W0_mask[2];
  assign mem_152_3_R0_addr = R0_addr[25:0];
  assign mem_152_3_R0_clk = R0_clk;
  assign mem_152_3_R0_en = R0_en & R0_addr_sel == 8'h98;
  assign mem_152_3_W0_addr = W0_addr[25:0];
  assign mem_152_3_W0_clk = W0_clk;
  assign mem_152_3_W0_data = W0_data[31:24];
  assign mem_152_3_W0_en = W0_en & W0_addr_sel == 8'h98;
  assign mem_152_3_W0_mask = W0_mask[3];
  assign mem_152_4_R0_addr = R0_addr[25:0];
  assign mem_152_4_R0_clk = R0_clk;
  assign mem_152_4_R0_en = R0_en & R0_addr_sel == 8'h98;
  assign mem_152_4_W0_addr = W0_addr[25:0];
  assign mem_152_4_W0_clk = W0_clk;
  assign mem_152_4_W0_data = W0_data[39:32];
  assign mem_152_4_W0_en = W0_en & W0_addr_sel == 8'h98;
  assign mem_152_4_W0_mask = W0_mask[4];
  assign mem_152_5_R0_addr = R0_addr[25:0];
  assign mem_152_5_R0_clk = R0_clk;
  assign mem_152_5_R0_en = R0_en & R0_addr_sel == 8'h98;
  assign mem_152_5_W0_addr = W0_addr[25:0];
  assign mem_152_5_W0_clk = W0_clk;
  assign mem_152_5_W0_data = W0_data[47:40];
  assign mem_152_5_W0_en = W0_en & W0_addr_sel == 8'h98;
  assign mem_152_5_W0_mask = W0_mask[5];
  assign mem_152_6_R0_addr = R0_addr[25:0];
  assign mem_152_6_R0_clk = R0_clk;
  assign mem_152_6_R0_en = R0_en & R0_addr_sel == 8'h98;
  assign mem_152_6_W0_addr = W0_addr[25:0];
  assign mem_152_6_W0_clk = W0_clk;
  assign mem_152_6_W0_data = W0_data[55:48];
  assign mem_152_6_W0_en = W0_en & W0_addr_sel == 8'h98;
  assign mem_152_6_W0_mask = W0_mask[6];
  assign mem_152_7_R0_addr = R0_addr[25:0];
  assign mem_152_7_R0_clk = R0_clk;
  assign mem_152_7_R0_en = R0_en & R0_addr_sel == 8'h98;
  assign mem_152_7_W0_addr = W0_addr[25:0];
  assign mem_152_7_W0_clk = W0_clk;
  assign mem_152_7_W0_data = W0_data[63:56];
  assign mem_152_7_W0_en = W0_en & W0_addr_sel == 8'h98;
  assign mem_152_7_W0_mask = W0_mask[7];
  assign mem_153_0_R0_addr = R0_addr[25:0];
  assign mem_153_0_R0_clk = R0_clk;
  assign mem_153_0_R0_en = R0_en & R0_addr_sel == 8'h99;
  assign mem_153_0_W0_addr = W0_addr[25:0];
  assign mem_153_0_W0_clk = W0_clk;
  assign mem_153_0_W0_data = W0_data[7:0];
  assign mem_153_0_W0_en = W0_en & W0_addr_sel == 8'h99;
  assign mem_153_0_W0_mask = W0_mask[0];
  assign mem_153_1_R0_addr = R0_addr[25:0];
  assign mem_153_1_R0_clk = R0_clk;
  assign mem_153_1_R0_en = R0_en & R0_addr_sel == 8'h99;
  assign mem_153_1_W0_addr = W0_addr[25:0];
  assign mem_153_1_W0_clk = W0_clk;
  assign mem_153_1_W0_data = W0_data[15:8];
  assign mem_153_1_W0_en = W0_en & W0_addr_sel == 8'h99;
  assign mem_153_1_W0_mask = W0_mask[1];
  assign mem_153_2_R0_addr = R0_addr[25:0];
  assign mem_153_2_R0_clk = R0_clk;
  assign mem_153_2_R0_en = R0_en & R0_addr_sel == 8'h99;
  assign mem_153_2_W0_addr = W0_addr[25:0];
  assign mem_153_2_W0_clk = W0_clk;
  assign mem_153_2_W0_data = W0_data[23:16];
  assign mem_153_2_W0_en = W0_en & W0_addr_sel == 8'h99;
  assign mem_153_2_W0_mask = W0_mask[2];
  assign mem_153_3_R0_addr = R0_addr[25:0];
  assign mem_153_3_R0_clk = R0_clk;
  assign mem_153_3_R0_en = R0_en & R0_addr_sel == 8'h99;
  assign mem_153_3_W0_addr = W0_addr[25:0];
  assign mem_153_3_W0_clk = W0_clk;
  assign mem_153_3_W0_data = W0_data[31:24];
  assign mem_153_3_W0_en = W0_en & W0_addr_sel == 8'h99;
  assign mem_153_3_W0_mask = W0_mask[3];
  assign mem_153_4_R0_addr = R0_addr[25:0];
  assign mem_153_4_R0_clk = R0_clk;
  assign mem_153_4_R0_en = R0_en & R0_addr_sel == 8'h99;
  assign mem_153_4_W0_addr = W0_addr[25:0];
  assign mem_153_4_W0_clk = W0_clk;
  assign mem_153_4_W0_data = W0_data[39:32];
  assign mem_153_4_W0_en = W0_en & W0_addr_sel == 8'h99;
  assign mem_153_4_W0_mask = W0_mask[4];
  assign mem_153_5_R0_addr = R0_addr[25:0];
  assign mem_153_5_R0_clk = R0_clk;
  assign mem_153_5_R0_en = R0_en & R0_addr_sel == 8'h99;
  assign mem_153_5_W0_addr = W0_addr[25:0];
  assign mem_153_5_W0_clk = W0_clk;
  assign mem_153_5_W0_data = W0_data[47:40];
  assign mem_153_5_W0_en = W0_en & W0_addr_sel == 8'h99;
  assign mem_153_5_W0_mask = W0_mask[5];
  assign mem_153_6_R0_addr = R0_addr[25:0];
  assign mem_153_6_R0_clk = R0_clk;
  assign mem_153_6_R0_en = R0_en & R0_addr_sel == 8'h99;
  assign mem_153_6_W0_addr = W0_addr[25:0];
  assign mem_153_6_W0_clk = W0_clk;
  assign mem_153_6_W0_data = W0_data[55:48];
  assign mem_153_6_W0_en = W0_en & W0_addr_sel == 8'h99;
  assign mem_153_6_W0_mask = W0_mask[6];
  assign mem_153_7_R0_addr = R0_addr[25:0];
  assign mem_153_7_R0_clk = R0_clk;
  assign mem_153_7_R0_en = R0_en & R0_addr_sel == 8'h99;
  assign mem_153_7_W0_addr = W0_addr[25:0];
  assign mem_153_7_W0_clk = W0_clk;
  assign mem_153_7_W0_data = W0_data[63:56];
  assign mem_153_7_W0_en = W0_en & W0_addr_sel == 8'h99;
  assign mem_153_7_W0_mask = W0_mask[7];
  assign mem_154_0_R0_addr = R0_addr[25:0];
  assign mem_154_0_R0_clk = R0_clk;
  assign mem_154_0_R0_en = R0_en & R0_addr_sel == 8'h9a;
  assign mem_154_0_W0_addr = W0_addr[25:0];
  assign mem_154_0_W0_clk = W0_clk;
  assign mem_154_0_W0_data = W0_data[7:0];
  assign mem_154_0_W0_en = W0_en & W0_addr_sel == 8'h9a;
  assign mem_154_0_W0_mask = W0_mask[0];
  assign mem_154_1_R0_addr = R0_addr[25:0];
  assign mem_154_1_R0_clk = R0_clk;
  assign mem_154_1_R0_en = R0_en & R0_addr_sel == 8'h9a;
  assign mem_154_1_W0_addr = W0_addr[25:0];
  assign mem_154_1_W0_clk = W0_clk;
  assign mem_154_1_W0_data = W0_data[15:8];
  assign mem_154_1_W0_en = W0_en & W0_addr_sel == 8'h9a;
  assign mem_154_1_W0_mask = W0_mask[1];
  assign mem_154_2_R0_addr = R0_addr[25:0];
  assign mem_154_2_R0_clk = R0_clk;
  assign mem_154_2_R0_en = R0_en & R0_addr_sel == 8'h9a;
  assign mem_154_2_W0_addr = W0_addr[25:0];
  assign mem_154_2_W0_clk = W0_clk;
  assign mem_154_2_W0_data = W0_data[23:16];
  assign mem_154_2_W0_en = W0_en & W0_addr_sel == 8'h9a;
  assign mem_154_2_W0_mask = W0_mask[2];
  assign mem_154_3_R0_addr = R0_addr[25:0];
  assign mem_154_3_R0_clk = R0_clk;
  assign mem_154_3_R0_en = R0_en & R0_addr_sel == 8'h9a;
  assign mem_154_3_W0_addr = W0_addr[25:0];
  assign mem_154_3_W0_clk = W0_clk;
  assign mem_154_3_W0_data = W0_data[31:24];
  assign mem_154_3_W0_en = W0_en & W0_addr_sel == 8'h9a;
  assign mem_154_3_W0_mask = W0_mask[3];
  assign mem_154_4_R0_addr = R0_addr[25:0];
  assign mem_154_4_R0_clk = R0_clk;
  assign mem_154_4_R0_en = R0_en & R0_addr_sel == 8'h9a;
  assign mem_154_4_W0_addr = W0_addr[25:0];
  assign mem_154_4_W0_clk = W0_clk;
  assign mem_154_4_W0_data = W0_data[39:32];
  assign mem_154_4_W0_en = W0_en & W0_addr_sel == 8'h9a;
  assign mem_154_4_W0_mask = W0_mask[4];
  assign mem_154_5_R0_addr = R0_addr[25:0];
  assign mem_154_5_R0_clk = R0_clk;
  assign mem_154_5_R0_en = R0_en & R0_addr_sel == 8'h9a;
  assign mem_154_5_W0_addr = W0_addr[25:0];
  assign mem_154_5_W0_clk = W0_clk;
  assign mem_154_5_W0_data = W0_data[47:40];
  assign mem_154_5_W0_en = W0_en & W0_addr_sel == 8'h9a;
  assign mem_154_5_W0_mask = W0_mask[5];
  assign mem_154_6_R0_addr = R0_addr[25:0];
  assign mem_154_6_R0_clk = R0_clk;
  assign mem_154_6_R0_en = R0_en & R0_addr_sel == 8'h9a;
  assign mem_154_6_W0_addr = W0_addr[25:0];
  assign mem_154_6_W0_clk = W0_clk;
  assign mem_154_6_W0_data = W0_data[55:48];
  assign mem_154_6_W0_en = W0_en & W0_addr_sel == 8'h9a;
  assign mem_154_6_W0_mask = W0_mask[6];
  assign mem_154_7_R0_addr = R0_addr[25:0];
  assign mem_154_7_R0_clk = R0_clk;
  assign mem_154_7_R0_en = R0_en & R0_addr_sel == 8'h9a;
  assign mem_154_7_W0_addr = W0_addr[25:0];
  assign mem_154_7_W0_clk = W0_clk;
  assign mem_154_7_W0_data = W0_data[63:56];
  assign mem_154_7_W0_en = W0_en & W0_addr_sel == 8'h9a;
  assign mem_154_7_W0_mask = W0_mask[7];
  assign mem_155_0_R0_addr = R0_addr[25:0];
  assign mem_155_0_R0_clk = R0_clk;
  assign mem_155_0_R0_en = R0_en & R0_addr_sel == 8'h9b;
  assign mem_155_0_W0_addr = W0_addr[25:0];
  assign mem_155_0_W0_clk = W0_clk;
  assign mem_155_0_W0_data = W0_data[7:0];
  assign mem_155_0_W0_en = W0_en & W0_addr_sel == 8'h9b;
  assign mem_155_0_W0_mask = W0_mask[0];
  assign mem_155_1_R0_addr = R0_addr[25:0];
  assign mem_155_1_R0_clk = R0_clk;
  assign mem_155_1_R0_en = R0_en & R0_addr_sel == 8'h9b;
  assign mem_155_1_W0_addr = W0_addr[25:0];
  assign mem_155_1_W0_clk = W0_clk;
  assign mem_155_1_W0_data = W0_data[15:8];
  assign mem_155_1_W0_en = W0_en & W0_addr_sel == 8'h9b;
  assign mem_155_1_W0_mask = W0_mask[1];
  assign mem_155_2_R0_addr = R0_addr[25:0];
  assign mem_155_2_R0_clk = R0_clk;
  assign mem_155_2_R0_en = R0_en & R0_addr_sel == 8'h9b;
  assign mem_155_2_W0_addr = W0_addr[25:0];
  assign mem_155_2_W0_clk = W0_clk;
  assign mem_155_2_W0_data = W0_data[23:16];
  assign mem_155_2_W0_en = W0_en & W0_addr_sel == 8'h9b;
  assign mem_155_2_W0_mask = W0_mask[2];
  assign mem_155_3_R0_addr = R0_addr[25:0];
  assign mem_155_3_R0_clk = R0_clk;
  assign mem_155_3_R0_en = R0_en & R0_addr_sel == 8'h9b;
  assign mem_155_3_W0_addr = W0_addr[25:0];
  assign mem_155_3_W0_clk = W0_clk;
  assign mem_155_3_W0_data = W0_data[31:24];
  assign mem_155_3_W0_en = W0_en & W0_addr_sel == 8'h9b;
  assign mem_155_3_W0_mask = W0_mask[3];
  assign mem_155_4_R0_addr = R0_addr[25:0];
  assign mem_155_4_R0_clk = R0_clk;
  assign mem_155_4_R0_en = R0_en & R0_addr_sel == 8'h9b;
  assign mem_155_4_W0_addr = W0_addr[25:0];
  assign mem_155_4_W0_clk = W0_clk;
  assign mem_155_4_W0_data = W0_data[39:32];
  assign mem_155_4_W0_en = W0_en & W0_addr_sel == 8'h9b;
  assign mem_155_4_W0_mask = W0_mask[4];
  assign mem_155_5_R0_addr = R0_addr[25:0];
  assign mem_155_5_R0_clk = R0_clk;
  assign mem_155_5_R0_en = R0_en & R0_addr_sel == 8'h9b;
  assign mem_155_5_W0_addr = W0_addr[25:0];
  assign mem_155_5_W0_clk = W0_clk;
  assign mem_155_5_W0_data = W0_data[47:40];
  assign mem_155_5_W0_en = W0_en & W0_addr_sel == 8'h9b;
  assign mem_155_5_W0_mask = W0_mask[5];
  assign mem_155_6_R0_addr = R0_addr[25:0];
  assign mem_155_6_R0_clk = R0_clk;
  assign mem_155_6_R0_en = R0_en & R0_addr_sel == 8'h9b;
  assign mem_155_6_W0_addr = W0_addr[25:0];
  assign mem_155_6_W0_clk = W0_clk;
  assign mem_155_6_W0_data = W0_data[55:48];
  assign mem_155_6_W0_en = W0_en & W0_addr_sel == 8'h9b;
  assign mem_155_6_W0_mask = W0_mask[6];
  assign mem_155_7_R0_addr = R0_addr[25:0];
  assign mem_155_7_R0_clk = R0_clk;
  assign mem_155_7_R0_en = R0_en & R0_addr_sel == 8'h9b;
  assign mem_155_7_W0_addr = W0_addr[25:0];
  assign mem_155_7_W0_clk = W0_clk;
  assign mem_155_7_W0_data = W0_data[63:56];
  assign mem_155_7_W0_en = W0_en & W0_addr_sel == 8'h9b;
  assign mem_155_7_W0_mask = W0_mask[7];
  assign mem_156_0_R0_addr = R0_addr[25:0];
  assign mem_156_0_R0_clk = R0_clk;
  assign mem_156_0_R0_en = R0_en & R0_addr_sel == 8'h9c;
  assign mem_156_0_W0_addr = W0_addr[25:0];
  assign mem_156_0_W0_clk = W0_clk;
  assign mem_156_0_W0_data = W0_data[7:0];
  assign mem_156_0_W0_en = W0_en & W0_addr_sel == 8'h9c;
  assign mem_156_0_W0_mask = W0_mask[0];
  assign mem_156_1_R0_addr = R0_addr[25:0];
  assign mem_156_1_R0_clk = R0_clk;
  assign mem_156_1_R0_en = R0_en & R0_addr_sel == 8'h9c;
  assign mem_156_1_W0_addr = W0_addr[25:0];
  assign mem_156_1_W0_clk = W0_clk;
  assign mem_156_1_W0_data = W0_data[15:8];
  assign mem_156_1_W0_en = W0_en & W0_addr_sel == 8'h9c;
  assign mem_156_1_W0_mask = W0_mask[1];
  assign mem_156_2_R0_addr = R0_addr[25:0];
  assign mem_156_2_R0_clk = R0_clk;
  assign mem_156_2_R0_en = R0_en & R0_addr_sel == 8'h9c;
  assign mem_156_2_W0_addr = W0_addr[25:0];
  assign mem_156_2_W0_clk = W0_clk;
  assign mem_156_2_W0_data = W0_data[23:16];
  assign mem_156_2_W0_en = W0_en & W0_addr_sel == 8'h9c;
  assign mem_156_2_W0_mask = W0_mask[2];
  assign mem_156_3_R0_addr = R0_addr[25:0];
  assign mem_156_3_R0_clk = R0_clk;
  assign mem_156_3_R0_en = R0_en & R0_addr_sel == 8'h9c;
  assign mem_156_3_W0_addr = W0_addr[25:0];
  assign mem_156_3_W0_clk = W0_clk;
  assign mem_156_3_W0_data = W0_data[31:24];
  assign mem_156_3_W0_en = W0_en & W0_addr_sel == 8'h9c;
  assign mem_156_3_W0_mask = W0_mask[3];
  assign mem_156_4_R0_addr = R0_addr[25:0];
  assign mem_156_4_R0_clk = R0_clk;
  assign mem_156_4_R0_en = R0_en & R0_addr_sel == 8'h9c;
  assign mem_156_4_W0_addr = W0_addr[25:0];
  assign mem_156_4_W0_clk = W0_clk;
  assign mem_156_4_W0_data = W0_data[39:32];
  assign mem_156_4_W0_en = W0_en & W0_addr_sel == 8'h9c;
  assign mem_156_4_W0_mask = W0_mask[4];
  assign mem_156_5_R0_addr = R0_addr[25:0];
  assign mem_156_5_R0_clk = R0_clk;
  assign mem_156_5_R0_en = R0_en & R0_addr_sel == 8'h9c;
  assign mem_156_5_W0_addr = W0_addr[25:0];
  assign mem_156_5_W0_clk = W0_clk;
  assign mem_156_5_W0_data = W0_data[47:40];
  assign mem_156_5_W0_en = W0_en & W0_addr_sel == 8'h9c;
  assign mem_156_5_W0_mask = W0_mask[5];
  assign mem_156_6_R0_addr = R0_addr[25:0];
  assign mem_156_6_R0_clk = R0_clk;
  assign mem_156_6_R0_en = R0_en & R0_addr_sel == 8'h9c;
  assign mem_156_6_W0_addr = W0_addr[25:0];
  assign mem_156_6_W0_clk = W0_clk;
  assign mem_156_6_W0_data = W0_data[55:48];
  assign mem_156_6_W0_en = W0_en & W0_addr_sel == 8'h9c;
  assign mem_156_6_W0_mask = W0_mask[6];
  assign mem_156_7_R0_addr = R0_addr[25:0];
  assign mem_156_7_R0_clk = R0_clk;
  assign mem_156_7_R0_en = R0_en & R0_addr_sel == 8'h9c;
  assign mem_156_7_W0_addr = W0_addr[25:0];
  assign mem_156_7_W0_clk = W0_clk;
  assign mem_156_7_W0_data = W0_data[63:56];
  assign mem_156_7_W0_en = W0_en & W0_addr_sel == 8'h9c;
  assign mem_156_7_W0_mask = W0_mask[7];
  assign mem_157_0_R0_addr = R0_addr[25:0];
  assign mem_157_0_R0_clk = R0_clk;
  assign mem_157_0_R0_en = R0_en & R0_addr_sel == 8'h9d;
  assign mem_157_0_W0_addr = W0_addr[25:0];
  assign mem_157_0_W0_clk = W0_clk;
  assign mem_157_0_W0_data = W0_data[7:0];
  assign mem_157_0_W0_en = W0_en & W0_addr_sel == 8'h9d;
  assign mem_157_0_W0_mask = W0_mask[0];
  assign mem_157_1_R0_addr = R0_addr[25:0];
  assign mem_157_1_R0_clk = R0_clk;
  assign mem_157_1_R0_en = R0_en & R0_addr_sel == 8'h9d;
  assign mem_157_1_W0_addr = W0_addr[25:0];
  assign mem_157_1_W0_clk = W0_clk;
  assign mem_157_1_W0_data = W0_data[15:8];
  assign mem_157_1_W0_en = W0_en & W0_addr_sel == 8'h9d;
  assign mem_157_1_W0_mask = W0_mask[1];
  assign mem_157_2_R0_addr = R0_addr[25:0];
  assign mem_157_2_R0_clk = R0_clk;
  assign mem_157_2_R0_en = R0_en & R0_addr_sel == 8'h9d;
  assign mem_157_2_W0_addr = W0_addr[25:0];
  assign mem_157_2_W0_clk = W0_clk;
  assign mem_157_2_W0_data = W0_data[23:16];
  assign mem_157_2_W0_en = W0_en & W0_addr_sel == 8'h9d;
  assign mem_157_2_W0_mask = W0_mask[2];
  assign mem_157_3_R0_addr = R0_addr[25:0];
  assign mem_157_3_R0_clk = R0_clk;
  assign mem_157_3_R0_en = R0_en & R0_addr_sel == 8'h9d;
  assign mem_157_3_W0_addr = W0_addr[25:0];
  assign mem_157_3_W0_clk = W0_clk;
  assign mem_157_3_W0_data = W0_data[31:24];
  assign mem_157_3_W0_en = W0_en & W0_addr_sel == 8'h9d;
  assign mem_157_3_W0_mask = W0_mask[3];
  assign mem_157_4_R0_addr = R0_addr[25:0];
  assign mem_157_4_R0_clk = R0_clk;
  assign mem_157_4_R0_en = R0_en & R0_addr_sel == 8'h9d;
  assign mem_157_4_W0_addr = W0_addr[25:0];
  assign mem_157_4_W0_clk = W0_clk;
  assign mem_157_4_W0_data = W0_data[39:32];
  assign mem_157_4_W0_en = W0_en & W0_addr_sel == 8'h9d;
  assign mem_157_4_W0_mask = W0_mask[4];
  assign mem_157_5_R0_addr = R0_addr[25:0];
  assign mem_157_5_R0_clk = R0_clk;
  assign mem_157_5_R0_en = R0_en & R0_addr_sel == 8'h9d;
  assign mem_157_5_W0_addr = W0_addr[25:0];
  assign mem_157_5_W0_clk = W0_clk;
  assign mem_157_5_W0_data = W0_data[47:40];
  assign mem_157_5_W0_en = W0_en & W0_addr_sel == 8'h9d;
  assign mem_157_5_W0_mask = W0_mask[5];
  assign mem_157_6_R0_addr = R0_addr[25:0];
  assign mem_157_6_R0_clk = R0_clk;
  assign mem_157_6_R0_en = R0_en & R0_addr_sel == 8'h9d;
  assign mem_157_6_W0_addr = W0_addr[25:0];
  assign mem_157_6_W0_clk = W0_clk;
  assign mem_157_6_W0_data = W0_data[55:48];
  assign mem_157_6_W0_en = W0_en & W0_addr_sel == 8'h9d;
  assign mem_157_6_W0_mask = W0_mask[6];
  assign mem_157_7_R0_addr = R0_addr[25:0];
  assign mem_157_7_R0_clk = R0_clk;
  assign mem_157_7_R0_en = R0_en & R0_addr_sel == 8'h9d;
  assign mem_157_7_W0_addr = W0_addr[25:0];
  assign mem_157_7_W0_clk = W0_clk;
  assign mem_157_7_W0_data = W0_data[63:56];
  assign mem_157_7_W0_en = W0_en & W0_addr_sel == 8'h9d;
  assign mem_157_7_W0_mask = W0_mask[7];
  assign mem_158_0_R0_addr = R0_addr[25:0];
  assign mem_158_0_R0_clk = R0_clk;
  assign mem_158_0_R0_en = R0_en & R0_addr_sel == 8'h9e;
  assign mem_158_0_W0_addr = W0_addr[25:0];
  assign mem_158_0_W0_clk = W0_clk;
  assign mem_158_0_W0_data = W0_data[7:0];
  assign mem_158_0_W0_en = W0_en & W0_addr_sel == 8'h9e;
  assign mem_158_0_W0_mask = W0_mask[0];
  assign mem_158_1_R0_addr = R0_addr[25:0];
  assign mem_158_1_R0_clk = R0_clk;
  assign mem_158_1_R0_en = R0_en & R0_addr_sel == 8'h9e;
  assign mem_158_1_W0_addr = W0_addr[25:0];
  assign mem_158_1_W0_clk = W0_clk;
  assign mem_158_1_W0_data = W0_data[15:8];
  assign mem_158_1_W0_en = W0_en & W0_addr_sel == 8'h9e;
  assign mem_158_1_W0_mask = W0_mask[1];
  assign mem_158_2_R0_addr = R0_addr[25:0];
  assign mem_158_2_R0_clk = R0_clk;
  assign mem_158_2_R0_en = R0_en & R0_addr_sel == 8'h9e;
  assign mem_158_2_W0_addr = W0_addr[25:0];
  assign mem_158_2_W0_clk = W0_clk;
  assign mem_158_2_W0_data = W0_data[23:16];
  assign mem_158_2_W0_en = W0_en & W0_addr_sel == 8'h9e;
  assign mem_158_2_W0_mask = W0_mask[2];
  assign mem_158_3_R0_addr = R0_addr[25:0];
  assign mem_158_3_R0_clk = R0_clk;
  assign mem_158_3_R0_en = R0_en & R0_addr_sel == 8'h9e;
  assign mem_158_3_W0_addr = W0_addr[25:0];
  assign mem_158_3_W0_clk = W0_clk;
  assign mem_158_3_W0_data = W0_data[31:24];
  assign mem_158_3_W0_en = W0_en & W0_addr_sel == 8'h9e;
  assign mem_158_3_W0_mask = W0_mask[3];
  assign mem_158_4_R0_addr = R0_addr[25:0];
  assign mem_158_4_R0_clk = R0_clk;
  assign mem_158_4_R0_en = R0_en & R0_addr_sel == 8'h9e;
  assign mem_158_4_W0_addr = W0_addr[25:0];
  assign mem_158_4_W0_clk = W0_clk;
  assign mem_158_4_W0_data = W0_data[39:32];
  assign mem_158_4_W0_en = W0_en & W0_addr_sel == 8'h9e;
  assign mem_158_4_W0_mask = W0_mask[4];
  assign mem_158_5_R0_addr = R0_addr[25:0];
  assign mem_158_5_R0_clk = R0_clk;
  assign mem_158_5_R0_en = R0_en & R0_addr_sel == 8'h9e;
  assign mem_158_5_W0_addr = W0_addr[25:0];
  assign mem_158_5_W0_clk = W0_clk;
  assign mem_158_5_W0_data = W0_data[47:40];
  assign mem_158_5_W0_en = W0_en & W0_addr_sel == 8'h9e;
  assign mem_158_5_W0_mask = W0_mask[5];
  assign mem_158_6_R0_addr = R0_addr[25:0];
  assign mem_158_6_R0_clk = R0_clk;
  assign mem_158_6_R0_en = R0_en & R0_addr_sel == 8'h9e;
  assign mem_158_6_W0_addr = W0_addr[25:0];
  assign mem_158_6_W0_clk = W0_clk;
  assign mem_158_6_W0_data = W0_data[55:48];
  assign mem_158_6_W0_en = W0_en & W0_addr_sel == 8'h9e;
  assign mem_158_6_W0_mask = W0_mask[6];
  assign mem_158_7_R0_addr = R0_addr[25:0];
  assign mem_158_7_R0_clk = R0_clk;
  assign mem_158_7_R0_en = R0_en & R0_addr_sel == 8'h9e;
  assign mem_158_7_W0_addr = W0_addr[25:0];
  assign mem_158_7_W0_clk = W0_clk;
  assign mem_158_7_W0_data = W0_data[63:56];
  assign mem_158_7_W0_en = W0_en & W0_addr_sel == 8'h9e;
  assign mem_158_7_W0_mask = W0_mask[7];
  assign mem_159_0_R0_addr = R0_addr[25:0];
  assign mem_159_0_R0_clk = R0_clk;
  assign mem_159_0_R0_en = R0_en & R0_addr_sel == 8'h9f;
  assign mem_159_0_W0_addr = W0_addr[25:0];
  assign mem_159_0_W0_clk = W0_clk;
  assign mem_159_0_W0_data = W0_data[7:0];
  assign mem_159_0_W0_en = W0_en & W0_addr_sel == 8'h9f;
  assign mem_159_0_W0_mask = W0_mask[0];
  assign mem_159_1_R0_addr = R0_addr[25:0];
  assign mem_159_1_R0_clk = R0_clk;
  assign mem_159_1_R0_en = R0_en & R0_addr_sel == 8'h9f;
  assign mem_159_1_W0_addr = W0_addr[25:0];
  assign mem_159_1_W0_clk = W0_clk;
  assign mem_159_1_W0_data = W0_data[15:8];
  assign mem_159_1_W0_en = W0_en & W0_addr_sel == 8'h9f;
  assign mem_159_1_W0_mask = W0_mask[1];
  assign mem_159_2_R0_addr = R0_addr[25:0];
  assign mem_159_2_R0_clk = R0_clk;
  assign mem_159_2_R0_en = R0_en & R0_addr_sel == 8'h9f;
  assign mem_159_2_W0_addr = W0_addr[25:0];
  assign mem_159_2_W0_clk = W0_clk;
  assign mem_159_2_W0_data = W0_data[23:16];
  assign mem_159_2_W0_en = W0_en & W0_addr_sel == 8'h9f;
  assign mem_159_2_W0_mask = W0_mask[2];
  assign mem_159_3_R0_addr = R0_addr[25:0];
  assign mem_159_3_R0_clk = R0_clk;
  assign mem_159_3_R0_en = R0_en & R0_addr_sel == 8'h9f;
  assign mem_159_3_W0_addr = W0_addr[25:0];
  assign mem_159_3_W0_clk = W0_clk;
  assign mem_159_3_W0_data = W0_data[31:24];
  assign mem_159_3_W0_en = W0_en & W0_addr_sel == 8'h9f;
  assign mem_159_3_W0_mask = W0_mask[3];
  assign mem_159_4_R0_addr = R0_addr[25:0];
  assign mem_159_4_R0_clk = R0_clk;
  assign mem_159_4_R0_en = R0_en & R0_addr_sel == 8'h9f;
  assign mem_159_4_W0_addr = W0_addr[25:0];
  assign mem_159_4_W0_clk = W0_clk;
  assign mem_159_4_W0_data = W0_data[39:32];
  assign mem_159_4_W0_en = W0_en & W0_addr_sel == 8'h9f;
  assign mem_159_4_W0_mask = W0_mask[4];
  assign mem_159_5_R0_addr = R0_addr[25:0];
  assign mem_159_5_R0_clk = R0_clk;
  assign mem_159_5_R0_en = R0_en & R0_addr_sel == 8'h9f;
  assign mem_159_5_W0_addr = W0_addr[25:0];
  assign mem_159_5_W0_clk = W0_clk;
  assign mem_159_5_W0_data = W0_data[47:40];
  assign mem_159_5_W0_en = W0_en & W0_addr_sel == 8'h9f;
  assign mem_159_5_W0_mask = W0_mask[5];
  assign mem_159_6_R0_addr = R0_addr[25:0];
  assign mem_159_6_R0_clk = R0_clk;
  assign mem_159_6_R0_en = R0_en & R0_addr_sel == 8'h9f;
  assign mem_159_6_W0_addr = W0_addr[25:0];
  assign mem_159_6_W0_clk = W0_clk;
  assign mem_159_6_W0_data = W0_data[55:48];
  assign mem_159_6_W0_en = W0_en & W0_addr_sel == 8'h9f;
  assign mem_159_6_W0_mask = W0_mask[6];
  assign mem_159_7_R0_addr = R0_addr[25:0];
  assign mem_159_7_R0_clk = R0_clk;
  assign mem_159_7_R0_en = R0_en & R0_addr_sel == 8'h9f;
  assign mem_159_7_W0_addr = W0_addr[25:0];
  assign mem_159_7_W0_clk = W0_clk;
  assign mem_159_7_W0_data = W0_data[63:56];
  assign mem_159_7_W0_en = W0_en & W0_addr_sel == 8'h9f;
  assign mem_159_7_W0_mask = W0_mask[7];
  assign mem_160_0_R0_addr = R0_addr[25:0];
  assign mem_160_0_R0_clk = R0_clk;
  assign mem_160_0_R0_en = R0_en & R0_addr_sel == 8'ha0;
  assign mem_160_0_W0_addr = W0_addr[25:0];
  assign mem_160_0_W0_clk = W0_clk;
  assign mem_160_0_W0_data = W0_data[7:0];
  assign mem_160_0_W0_en = W0_en & W0_addr_sel == 8'ha0;
  assign mem_160_0_W0_mask = W0_mask[0];
  assign mem_160_1_R0_addr = R0_addr[25:0];
  assign mem_160_1_R0_clk = R0_clk;
  assign mem_160_1_R0_en = R0_en & R0_addr_sel == 8'ha0;
  assign mem_160_1_W0_addr = W0_addr[25:0];
  assign mem_160_1_W0_clk = W0_clk;
  assign mem_160_1_W0_data = W0_data[15:8];
  assign mem_160_1_W0_en = W0_en & W0_addr_sel == 8'ha0;
  assign mem_160_1_W0_mask = W0_mask[1];
  assign mem_160_2_R0_addr = R0_addr[25:0];
  assign mem_160_2_R0_clk = R0_clk;
  assign mem_160_2_R0_en = R0_en & R0_addr_sel == 8'ha0;
  assign mem_160_2_W0_addr = W0_addr[25:0];
  assign mem_160_2_W0_clk = W0_clk;
  assign mem_160_2_W0_data = W0_data[23:16];
  assign mem_160_2_W0_en = W0_en & W0_addr_sel == 8'ha0;
  assign mem_160_2_W0_mask = W0_mask[2];
  assign mem_160_3_R0_addr = R0_addr[25:0];
  assign mem_160_3_R0_clk = R0_clk;
  assign mem_160_3_R0_en = R0_en & R0_addr_sel == 8'ha0;
  assign mem_160_3_W0_addr = W0_addr[25:0];
  assign mem_160_3_W0_clk = W0_clk;
  assign mem_160_3_W0_data = W0_data[31:24];
  assign mem_160_3_W0_en = W0_en & W0_addr_sel == 8'ha0;
  assign mem_160_3_W0_mask = W0_mask[3];
  assign mem_160_4_R0_addr = R0_addr[25:0];
  assign mem_160_4_R0_clk = R0_clk;
  assign mem_160_4_R0_en = R0_en & R0_addr_sel == 8'ha0;
  assign mem_160_4_W0_addr = W0_addr[25:0];
  assign mem_160_4_W0_clk = W0_clk;
  assign mem_160_4_W0_data = W0_data[39:32];
  assign mem_160_4_W0_en = W0_en & W0_addr_sel == 8'ha0;
  assign mem_160_4_W0_mask = W0_mask[4];
  assign mem_160_5_R0_addr = R0_addr[25:0];
  assign mem_160_5_R0_clk = R0_clk;
  assign mem_160_5_R0_en = R0_en & R0_addr_sel == 8'ha0;
  assign mem_160_5_W0_addr = W0_addr[25:0];
  assign mem_160_5_W0_clk = W0_clk;
  assign mem_160_5_W0_data = W0_data[47:40];
  assign mem_160_5_W0_en = W0_en & W0_addr_sel == 8'ha0;
  assign mem_160_5_W0_mask = W0_mask[5];
  assign mem_160_6_R0_addr = R0_addr[25:0];
  assign mem_160_6_R0_clk = R0_clk;
  assign mem_160_6_R0_en = R0_en & R0_addr_sel == 8'ha0;
  assign mem_160_6_W0_addr = W0_addr[25:0];
  assign mem_160_6_W0_clk = W0_clk;
  assign mem_160_6_W0_data = W0_data[55:48];
  assign mem_160_6_W0_en = W0_en & W0_addr_sel == 8'ha0;
  assign mem_160_6_W0_mask = W0_mask[6];
  assign mem_160_7_R0_addr = R0_addr[25:0];
  assign mem_160_7_R0_clk = R0_clk;
  assign mem_160_7_R0_en = R0_en & R0_addr_sel == 8'ha0;
  assign mem_160_7_W0_addr = W0_addr[25:0];
  assign mem_160_7_W0_clk = W0_clk;
  assign mem_160_7_W0_data = W0_data[63:56];
  assign mem_160_7_W0_en = W0_en & W0_addr_sel == 8'ha0;
  assign mem_160_7_W0_mask = W0_mask[7];
  assign mem_161_0_R0_addr = R0_addr[25:0];
  assign mem_161_0_R0_clk = R0_clk;
  assign mem_161_0_R0_en = R0_en & R0_addr_sel == 8'ha1;
  assign mem_161_0_W0_addr = W0_addr[25:0];
  assign mem_161_0_W0_clk = W0_clk;
  assign mem_161_0_W0_data = W0_data[7:0];
  assign mem_161_0_W0_en = W0_en & W0_addr_sel == 8'ha1;
  assign mem_161_0_W0_mask = W0_mask[0];
  assign mem_161_1_R0_addr = R0_addr[25:0];
  assign mem_161_1_R0_clk = R0_clk;
  assign mem_161_1_R0_en = R0_en & R0_addr_sel == 8'ha1;
  assign mem_161_1_W0_addr = W0_addr[25:0];
  assign mem_161_1_W0_clk = W0_clk;
  assign mem_161_1_W0_data = W0_data[15:8];
  assign mem_161_1_W0_en = W0_en & W0_addr_sel == 8'ha1;
  assign mem_161_1_W0_mask = W0_mask[1];
  assign mem_161_2_R0_addr = R0_addr[25:0];
  assign mem_161_2_R0_clk = R0_clk;
  assign mem_161_2_R0_en = R0_en & R0_addr_sel == 8'ha1;
  assign mem_161_2_W0_addr = W0_addr[25:0];
  assign mem_161_2_W0_clk = W0_clk;
  assign mem_161_2_W0_data = W0_data[23:16];
  assign mem_161_2_W0_en = W0_en & W0_addr_sel == 8'ha1;
  assign mem_161_2_W0_mask = W0_mask[2];
  assign mem_161_3_R0_addr = R0_addr[25:0];
  assign mem_161_3_R0_clk = R0_clk;
  assign mem_161_3_R0_en = R0_en & R0_addr_sel == 8'ha1;
  assign mem_161_3_W0_addr = W0_addr[25:0];
  assign mem_161_3_W0_clk = W0_clk;
  assign mem_161_3_W0_data = W0_data[31:24];
  assign mem_161_3_W0_en = W0_en & W0_addr_sel == 8'ha1;
  assign mem_161_3_W0_mask = W0_mask[3];
  assign mem_161_4_R0_addr = R0_addr[25:0];
  assign mem_161_4_R0_clk = R0_clk;
  assign mem_161_4_R0_en = R0_en & R0_addr_sel == 8'ha1;
  assign mem_161_4_W0_addr = W0_addr[25:0];
  assign mem_161_4_W0_clk = W0_clk;
  assign mem_161_4_W0_data = W0_data[39:32];
  assign mem_161_4_W0_en = W0_en & W0_addr_sel == 8'ha1;
  assign mem_161_4_W0_mask = W0_mask[4];
  assign mem_161_5_R0_addr = R0_addr[25:0];
  assign mem_161_5_R0_clk = R0_clk;
  assign mem_161_5_R0_en = R0_en & R0_addr_sel == 8'ha1;
  assign mem_161_5_W0_addr = W0_addr[25:0];
  assign mem_161_5_W0_clk = W0_clk;
  assign mem_161_5_W0_data = W0_data[47:40];
  assign mem_161_5_W0_en = W0_en & W0_addr_sel == 8'ha1;
  assign mem_161_5_W0_mask = W0_mask[5];
  assign mem_161_6_R0_addr = R0_addr[25:0];
  assign mem_161_6_R0_clk = R0_clk;
  assign mem_161_6_R0_en = R0_en & R0_addr_sel == 8'ha1;
  assign mem_161_6_W0_addr = W0_addr[25:0];
  assign mem_161_6_W0_clk = W0_clk;
  assign mem_161_6_W0_data = W0_data[55:48];
  assign mem_161_6_W0_en = W0_en & W0_addr_sel == 8'ha1;
  assign mem_161_6_W0_mask = W0_mask[6];
  assign mem_161_7_R0_addr = R0_addr[25:0];
  assign mem_161_7_R0_clk = R0_clk;
  assign mem_161_7_R0_en = R0_en & R0_addr_sel == 8'ha1;
  assign mem_161_7_W0_addr = W0_addr[25:0];
  assign mem_161_7_W0_clk = W0_clk;
  assign mem_161_7_W0_data = W0_data[63:56];
  assign mem_161_7_W0_en = W0_en & W0_addr_sel == 8'ha1;
  assign mem_161_7_W0_mask = W0_mask[7];
  assign mem_162_0_R0_addr = R0_addr[25:0];
  assign mem_162_0_R0_clk = R0_clk;
  assign mem_162_0_R0_en = R0_en & R0_addr_sel == 8'ha2;
  assign mem_162_0_W0_addr = W0_addr[25:0];
  assign mem_162_0_W0_clk = W0_clk;
  assign mem_162_0_W0_data = W0_data[7:0];
  assign mem_162_0_W0_en = W0_en & W0_addr_sel == 8'ha2;
  assign mem_162_0_W0_mask = W0_mask[0];
  assign mem_162_1_R0_addr = R0_addr[25:0];
  assign mem_162_1_R0_clk = R0_clk;
  assign mem_162_1_R0_en = R0_en & R0_addr_sel == 8'ha2;
  assign mem_162_1_W0_addr = W0_addr[25:0];
  assign mem_162_1_W0_clk = W0_clk;
  assign mem_162_1_W0_data = W0_data[15:8];
  assign mem_162_1_W0_en = W0_en & W0_addr_sel == 8'ha2;
  assign mem_162_1_W0_mask = W0_mask[1];
  assign mem_162_2_R0_addr = R0_addr[25:0];
  assign mem_162_2_R0_clk = R0_clk;
  assign mem_162_2_R0_en = R0_en & R0_addr_sel == 8'ha2;
  assign mem_162_2_W0_addr = W0_addr[25:0];
  assign mem_162_2_W0_clk = W0_clk;
  assign mem_162_2_W0_data = W0_data[23:16];
  assign mem_162_2_W0_en = W0_en & W0_addr_sel == 8'ha2;
  assign mem_162_2_W0_mask = W0_mask[2];
  assign mem_162_3_R0_addr = R0_addr[25:0];
  assign mem_162_3_R0_clk = R0_clk;
  assign mem_162_3_R0_en = R0_en & R0_addr_sel == 8'ha2;
  assign mem_162_3_W0_addr = W0_addr[25:0];
  assign mem_162_3_W0_clk = W0_clk;
  assign mem_162_3_W0_data = W0_data[31:24];
  assign mem_162_3_W0_en = W0_en & W0_addr_sel == 8'ha2;
  assign mem_162_3_W0_mask = W0_mask[3];
  assign mem_162_4_R0_addr = R0_addr[25:0];
  assign mem_162_4_R0_clk = R0_clk;
  assign mem_162_4_R0_en = R0_en & R0_addr_sel == 8'ha2;
  assign mem_162_4_W0_addr = W0_addr[25:0];
  assign mem_162_4_W0_clk = W0_clk;
  assign mem_162_4_W0_data = W0_data[39:32];
  assign mem_162_4_W0_en = W0_en & W0_addr_sel == 8'ha2;
  assign mem_162_4_W0_mask = W0_mask[4];
  assign mem_162_5_R0_addr = R0_addr[25:0];
  assign mem_162_5_R0_clk = R0_clk;
  assign mem_162_5_R0_en = R0_en & R0_addr_sel == 8'ha2;
  assign mem_162_5_W0_addr = W0_addr[25:0];
  assign mem_162_5_W0_clk = W0_clk;
  assign mem_162_5_W0_data = W0_data[47:40];
  assign mem_162_5_W0_en = W0_en & W0_addr_sel == 8'ha2;
  assign mem_162_5_W0_mask = W0_mask[5];
  assign mem_162_6_R0_addr = R0_addr[25:0];
  assign mem_162_6_R0_clk = R0_clk;
  assign mem_162_6_R0_en = R0_en & R0_addr_sel == 8'ha2;
  assign mem_162_6_W0_addr = W0_addr[25:0];
  assign mem_162_6_W0_clk = W0_clk;
  assign mem_162_6_W0_data = W0_data[55:48];
  assign mem_162_6_W0_en = W0_en & W0_addr_sel == 8'ha2;
  assign mem_162_6_W0_mask = W0_mask[6];
  assign mem_162_7_R0_addr = R0_addr[25:0];
  assign mem_162_7_R0_clk = R0_clk;
  assign mem_162_7_R0_en = R0_en & R0_addr_sel == 8'ha2;
  assign mem_162_7_W0_addr = W0_addr[25:0];
  assign mem_162_7_W0_clk = W0_clk;
  assign mem_162_7_W0_data = W0_data[63:56];
  assign mem_162_7_W0_en = W0_en & W0_addr_sel == 8'ha2;
  assign mem_162_7_W0_mask = W0_mask[7];
  assign mem_163_0_R0_addr = R0_addr[25:0];
  assign mem_163_0_R0_clk = R0_clk;
  assign mem_163_0_R0_en = R0_en & R0_addr_sel == 8'ha3;
  assign mem_163_0_W0_addr = W0_addr[25:0];
  assign mem_163_0_W0_clk = W0_clk;
  assign mem_163_0_W0_data = W0_data[7:0];
  assign mem_163_0_W0_en = W0_en & W0_addr_sel == 8'ha3;
  assign mem_163_0_W0_mask = W0_mask[0];
  assign mem_163_1_R0_addr = R0_addr[25:0];
  assign mem_163_1_R0_clk = R0_clk;
  assign mem_163_1_R0_en = R0_en & R0_addr_sel == 8'ha3;
  assign mem_163_1_W0_addr = W0_addr[25:0];
  assign mem_163_1_W0_clk = W0_clk;
  assign mem_163_1_W0_data = W0_data[15:8];
  assign mem_163_1_W0_en = W0_en & W0_addr_sel == 8'ha3;
  assign mem_163_1_W0_mask = W0_mask[1];
  assign mem_163_2_R0_addr = R0_addr[25:0];
  assign mem_163_2_R0_clk = R0_clk;
  assign mem_163_2_R0_en = R0_en & R0_addr_sel == 8'ha3;
  assign mem_163_2_W0_addr = W0_addr[25:0];
  assign mem_163_2_W0_clk = W0_clk;
  assign mem_163_2_W0_data = W0_data[23:16];
  assign mem_163_2_W0_en = W0_en & W0_addr_sel == 8'ha3;
  assign mem_163_2_W0_mask = W0_mask[2];
  assign mem_163_3_R0_addr = R0_addr[25:0];
  assign mem_163_3_R0_clk = R0_clk;
  assign mem_163_3_R0_en = R0_en & R0_addr_sel == 8'ha3;
  assign mem_163_3_W0_addr = W0_addr[25:0];
  assign mem_163_3_W0_clk = W0_clk;
  assign mem_163_3_W0_data = W0_data[31:24];
  assign mem_163_3_W0_en = W0_en & W0_addr_sel == 8'ha3;
  assign mem_163_3_W0_mask = W0_mask[3];
  assign mem_163_4_R0_addr = R0_addr[25:0];
  assign mem_163_4_R0_clk = R0_clk;
  assign mem_163_4_R0_en = R0_en & R0_addr_sel == 8'ha3;
  assign mem_163_4_W0_addr = W0_addr[25:0];
  assign mem_163_4_W0_clk = W0_clk;
  assign mem_163_4_W0_data = W0_data[39:32];
  assign mem_163_4_W0_en = W0_en & W0_addr_sel == 8'ha3;
  assign mem_163_4_W0_mask = W0_mask[4];
  assign mem_163_5_R0_addr = R0_addr[25:0];
  assign mem_163_5_R0_clk = R0_clk;
  assign mem_163_5_R0_en = R0_en & R0_addr_sel == 8'ha3;
  assign mem_163_5_W0_addr = W0_addr[25:0];
  assign mem_163_5_W0_clk = W0_clk;
  assign mem_163_5_W0_data = W0_data[47:40];
  assign mem_163_5_W0_en = W0_en & W0_addr_sel == 8'ha3;
  assign mem_163_5_W0_mask = W0_mask[5];
  assign mem_163_6_R0_addr = R0_addr[25:0];
  assign mem_163_6_R0_clk = R0_clk;
  assign mem_163_6_R0_en = R0_en & R0_addr_sel == 8'ha3;
  assign mem_163_6_W0_addr = W0_addr[25:0];
  assign mem_163_6_W0_clk = W0_clk;
  assign mem_163_6_W0_data = W0_data[55:48];
  assign mem_163_6_W0_en = W0_en & W0_addr_sel == 8'ha3;
  assign mem_163_6_W0_mask = W0_mask[6];
  assign mem_163_7_R0_addr = R0_addr[25:0];
  assign mem_163_7_R0_clk = R0_clk;
  assign mem_163_7_R0_en = R0_en & R0_addr_sel == 8'ha3;
  assign mem_163_7_W0_addr = W0_addr[25:0];
  assign mem_163_7_W0_clk = W0_clk;
  assign mem_163_7_W0_data = W0_data[63:56];
  assign mem_163_7_W0_en = W0_en & W0_addr_sel == 8'ha3;
  assign mem_163_7_W0_mask = W0_mask[7];
  assign mem_164_0_R0_addr = R0_addr[25:0];
  assign mem_164_0_R0_clk = R0_clk;
  assign mem_164_0_R0_en = R0_en & R0_addr_sel == 8'ha4;
  assign mem_164_0_W0_addr = W0_addr[25:0];
  assign mem_164_0_W0_clk = W0_clk;
  assign mem_164_0_W0_data = W0_data[7:0];
  assign mem_164_0_W0_en = W0_en & W0_addr_sel == 8'ha4;
  assign mem_164_0_W0_mask = W0_mask[0];
  assign mem_164_1_R0_addr = R0_addr[25:0];
  assign mem_164_1_R0_clk = R0_clk;
  assign mem_164_1_R0_en = R0_en & R0_addr_sel == 8'ha4;
  assign mem_164_1_W0_addr = W0_addr[25:0];
  assign mem_164_1_W0_clk = W0_clk;
  assign mem_164_1_W0_data = W0_data[15:8];
  assign mem_164_1_W0_en = W0_en & W0_addr_sel == 8'ha4;
  assign mem_164_1_W0_mask = W0_mask[1];
  assign mem_164_2_R0_addr = R0_addr[25:0];
  assign mem_164_2_R0_clk = R0_clk;
  assign mem_164_2_R0_en = R0_en & R0_addr_sel == 8'ha4;
  assign mem_164_2_W0_addr = W0_addr[25:0];
  assign mem_164_2_W0_clk = W0_clk;
  assign mem_164_2_W0_data = W0_data[23:16];
  assign mem_164_2_W0_en = W0_en & W0_addr_sel == 8'ha4;
  assign mem_164_2_W0_mask = W0_mask[2];
  assign mem_164_3_R0_addr = R0_addr[25:0];
  assign mem_164_3_R0_clk = R0_clk;
  assign mem_164_3_R0_en = R0_en & R0_addr_sel == 8'ha4;
  assign mem_164_3_W0_addr = W0_addr[25:0];
  assign mem_164_3_W0_clk = W0_clk;
  assign mem_164_3_W0_data = W0_data[31:24];
  assign mem_164_3_W0_en = W0_en & W0_addr_sel == 8'ha4;
  assign mem_164_3_W0_mask = W0_mask[3];
  assign mem_164_4_R0_addr = R0_addr[25:0];
  assign mem_164_4_R0_clk = R0_clk;
  assign mem_164_4_R0_en = R0_en & R0_addr_sel == 8'ha4;
  assign mem_164_4_W0_addr = W0_addr[25:0];
  assign mem_164_4_W0_clk = W0_clk;
  assign mem_164_4_W0_data = W0_data[39:32];
  assign mem_164_4_W0_en = W0_en & W0_addr_sel == 8'ha4;
  assign mem_164_4_W0_mask = W0_mask[4];
  assign mem_164_5_R0_addr = R0_addr[25:0];
  assign mem_164_5_R0_clk = R0_clk;
  assign mem_164_5_R0_en = R0_en & R0_addr_sel == 8'ha4;
  assign mem_164_5_W0_addr = W0_addr[25:0];
  assign mem_164_5_W0_clk = W0_clk;
  assign mem_164_5_W0_data = W0_data[47:40];
  assign mem_164_5_W0_en = W0_en & W0_addr_sel == 8'ha4;
  assign mem_164_5_W0_mask = W0_mask[5];
  assign mem_164_6_R0_addr = R0_addr[25:0];
  assign mem_164_6_R0_clk = R0_clk;
  assign mem_164_6_R0_en = R0_en & R0_addr_sel == 8'ha4;
  assign mem_164_6_W0_addr = W0_addr[25:0];
  assign mem_164_6_W0_clk = W0_clk;
  assign mem_164_6_W0_data = W0_data[55:48];
  assign mem_164_6_W0_en = W0_en & W0_addr_sel == 8'ha4;
  assign mem_164_6_W0_mask = W0_mask[6];
  assign mem_164_7_R0_addr = R0_addr[25:0];
  assign mem_164_7_R0_clk = R0_clk;
  assign mem_164_7_R0_en = R0_en & R0_addr_sel == 8'ha4;
  assign mem_164_7_W0_addr = W0_addr[25:0];
  assign mem_164_7_W0_clk = W0_clk;
  assign mem_164_7_W0_data = W0_data[63:56];
  assign mem_164_7_W0_en = W0_en & W0_addr_sel == 8'ha4;
  assign mem_164_7_W0_mask = W0_mask[7];
  assign mem_165_0_R0_addr = R0_addr[25:0];
  assign mem_165_0_R0_clk = R0_clk;
  assign mem_165_0_R0_en = R0_en & R0_addr_sel == 8'ha5;
  assign mem_165_0_W0_addr = W0_addr[25:0];
  assign mem_165_0_W0_clk = W0_clk;
  assign mem_165_0_W0_data = W0_data[7:0];
  assign mem_165_0_W0_en = W0_en & W0_addr_sel == 8'ha5;
  assign mem_165_0_W0_mask = W0_mask[0];
  assign mem_165_1_R0_addr = R0_addr[25:0];
  assign mem_165_1_R0_clk = R0_clk;
  assign mem_165_1_R0_en = R0_en & R0_addr_sel == 8'ha5;
  assign mem_165_1_W0_addr = W0_addr[25:0];
  assign mem_165_1_W0_clk = W0_clk;
  assign mem_165_1_W0_data = W0_data[15:8];
  assign mem_165_1_W0_en = W0_en & W0_addr_sel == 8'ha5;
  assign mem_165_1_W0_mask = W0_mask[1];
  assign mem_165_2_R0_addr = R0_addr[25:0];
  assign mem_165_2_R0_clk = R0_clk;
  assign mem_165_2_R0_en = R0_en & R0_addr_sel == 8'ha5;
  assign mem_165_2_W0_addr = W0_addr[25:0];
  assign mem_165_2_W0_clk = W0_clk;
  assign mem_165_2_W0_data = W0_data[23:16];
  assign mem_165_2_W0_en = W0_en & W0_addr_sel == 8'ha5;
  assign mem_165_2_W0_mask = W0_mask[2];
  assign mem_165_3_R0_addr = R0_addr[25:0];
  assign mem_165_3_R0_clk = R0_clk;
  assign mem_165_3_R0_en = R0_en & R0_addr_sel == 8'ha5;
  assign mem_165_3_W0_addr = W0_addr[25:0];
  assign mem_165_3_W0_clk = W0_clk;
  assign mem_165_3_W0_data = W0_data[31:24];
  assign mem_165_3_W0_en = W0_en & W0_addr_sel == 8'ha5;
  assign mem_165_3_W0_mask = W0_mask[3];
  assign mem_165_4_R0_addr = R0_addr[25:0];
  assign mem_165_4_R0_clk = R0_clk;
  assign mem_165_4_R0_en = R0_en & R0_addr_sel == 8'ha5;
  assign mem_165_4_W0_addr = W0_addr[25:0];
  assign mem_165_4_W0_clk = W0_clk;
  assign mem_165_4_W0_data = W0_data[39:32];
  assign mem_165_4_W0_en = W0_en & W0_addr_sel == 8'ha5;
  assign mem_165_4_W0_mask = W0_mask[4];
  assign mem_165_5_R0_addr = R0_addr[25:0];
  assign mem_165_5_R0_clk = R0_clk;
  assign mem_165_5_R0_en = R0_en & R0_addr_sel == 8'ha5;
  assign mem_165_5_W0_addr = W0_addr[25:0];
  assign mem_165_5_W0_clk = W0_clk;
  assign mem_165_5_W0_data = W0_data[47:40];
  assign mem_165_5_W0_en = W0_en & W0_addr_sel == 8'ha5;
  assign mem_165_5_W0_mask = W0_mask[5];
  assign mem_165_6_R0_addr = R0_addr[25:0];
  assign mem_165_6_R0_clk = R0_clk;
  assign mem_165_6_R0_en = R0_en & R0_addr_sel == 8'ha5;
  assign mem_165_6_W0_addr = W0_addr[25:0];
  assign mem_165_6_W0_clk = W0_clk;
  assign mem_165_6_W0_data = W0_data[55:48];
  assign mem_165_6_W0_en = W0_en & W0_addr_sel == 8'ha5;
  assign mem_165_6_W0_mask = W0_mask[6];
  assign mem_165_7_R0_addr = R0_addr[25:0];
  assign mem_165_7_R0_clk = R0_clk;
  assign mem_165_7_R0_en = R0_en & R0_addr_sel == 8'ha5;
  assign mem_165_7_W0_addr = W0_addr[25:0];
  assign mem_165_7_W0_clk = W0_clk;
  assign mem_165_7_W0_data = W0_data[63:56];
  assign mem_165_7_W0_en = W0_en & W0_addr_sel == 8'ha5;
  assign mem_165_7_W0_mask = W0_mask[7];
  assign mem_166_0_R0_addr = R0_addr[25:0];
  assign mem_166_0_R0_clk = R0_clk;
  assign mem_166_0_R0_en = R0_en & R0_addr_sel == 8'ha6;
  assign mem_166_0_W0_addr = W0_addr[25:0];
  assign mem_166_0_W0_clk = W0_clk;
  assign mem_166_0_W0_data = W0_data[7:0];
  assign mem_166_0_W0_en = W0_en & W0_addr_sel == 8'ha6;
  assign mem_166_0_W0_mask = W0_mask[0];
  assign mem_166_1_R0_addr = R0_addr[25:0];
  assign mem_166_1_R0_clk = R0_clk;
  assign mem_166_1_R0_en = R0_en & R0_addr_sel == 8'ha6;
  assign mem_166_1_W0_addr = W0_addr[25:0];
  assign mem_166_1_W0_clk = W0_clk;
  assign mem_166_1_W0_data = W0_data[15:8];
  assign mem_166_1_W0_en = W0_en & W0_addr_sel == 8'ha6;
  assign mem_166_1_W0_mask = W0_mask[1];
  assign mem_166_2_R0_addr = R0_addr[25:0];
  assign mem_166_2_R0_clk = R0_clk;
  assign mem_166_2_R0_en = R0_en & R0_addr_sel == 8'ha6;
  assign mem_166_2_W0_addr = W0_addr[25:0];
  assign mem_166_2_W0_clk = W0_clk;
  assign mem_166_2_W0_data = W0_data[23:16];
  assign mem_166_2_W0_en = W0_en & W0_addr_sel == 8'ha6;
  assign mem_166_2_W0_mask = W0_mask[2];
  assign mem_166_3_R0_addr = R0_addr[25:0];
  assign mem_166_3_R0_clk = R0_clk;
  assign mem_166_3_R0_en = R0_en & R0_addr_sel == 8'ha6;
  assign mem_166_3_W0_addr = W0_addr[25:0];
  assign mem_166_3_W0_clk = W0_clk;
  assign mem_166_3_W0_data = W0_data[31:24];
  assign mem_166_3_W0_en = W0_en & W0_addr_sel == 8'ha6;
  assign mem_166_3_W0_mask = W0_mask[3];
  assign mem_166_4_R0_addr = R0_addr[25:0];
  assign mem_166_4_R0_clk = R0_clk;
  assign mem_166_4_R0_en = R0_en & R0_addr_sel == 8'ha6;
  assign mem_166_4_W0_addr = W0_addr[25:0];
  assign mem_166_4_W0_clk = W0_clk;
  assign mem_166_4_W0_data = W0_data[39:32];
  assign mem_166_4_W0_en = W0_en & W0_addr_sel == 8'ha6;
  assign mem_166_4_W0_mask = W0_mask[4];
  assign mem_166_5_R0_addr = R0_addr[25:0];
  assign mem_166_5_R0_clk = R0_clk;
  assign mem_166_5_R0_en = R0_en & R0_addr_sel == 8'ha6;
  assign mem_166_5_W0_addr = W0_addr[25:0];
  assign mem_166_5_W0_clk = W0_clk;
  assign mem_166_5_W0_data = W0_data[47:40];
  assign mem_166_5_W0_en = W0_en & W0_addr_sel == 8'ha6;
  assign mem_166_5_W0_mask = W0_mask[5];
  assign mem_166_6_R0_addr = R0_addr[25:0];
  assign mem_166_6_R0_clk = R0_clk;
  assign mem_166_6_R0_en = R0_en & R0_addr_sel == 8'ha6;
  assign mem_166_6_W0_addr = W0_addr[25:0];
  assign mem_166_6_W0_clk = W0_clk;
  assign mem_166_6_W0_data = W0_data[55:48];
  assign mem_166_6_W0_en = W0_en & W0_addr_sel == 8'ha6;
  assign mem_166_6_W0_mask = W0_mask[6];
  assign mem_166_7_R0_addr = R0_addr[25:0];
  assign mem_166_7_R0_clk = R0_clk;
  assign mem_166_7_R0_en = R0_en & R0_addr_sel == 8'ha6;
  assign mem_166_7_W0_addr = W0_addr[25:0];
  assign mem_166_7_W0_clk = W0_clk;
  assign mem_166_7_W0_data = W0_data[63:56];
  assign mem_166_7_W0_en = W0_en & W0_addr_sel == 8'ha6;
  assign mem_166_7_W0_mask = W0_mask[7];
  assign mem_167_0_R0_addr = R0_addr[25:0];
  assign mem_167_0_R0_clk = R0_clk;
  assign mem_167_0_R0_en = R0_en & R0_addr_sel == 8'ha7;
  assign mem_167_0_W0_addr = W0_addr[25:0];
  assign mem_167_0_W0_clk = W0_clk;
  assign mem_167_0_W0_data = W0_data[7:0];
  assign mem_167_0_W0_en = W0_en & W0_addr_sel == 8'ha7;
  assign mem_167_0_W0_mask = W0_mask[0];
  assign mem_167_1_R0_addr = R0_addr[25:0];
  assign mem_167_1_R0_clk = R0_clk;
  assign mem_167_1_R0_en = R0_en & R0_addr_sel == 8'ha7;
  assign mem_167_1_W0_addr = W0_addr[25:0];
  assign mem_167_1_W0_clk = W0_clk;
  assign mem_167_1_W0_data = W0_data[15:8];
  assign mem_167_1_W0_en = W0_en & W0_addr_sel == 8'ha7;
  assign mem_167_1_W0_mask = W0_mask[1];
  assign mem_167_2_R0_addr = R0_addr[25:0];
  assign mem_167_2_R0_clk = R0_clk;
  assign mem_167_2_R0_en = R0_en & R0_addr_sel == 8'ha7;
  assign mem_167_2_W0_addr = W0_addr[25:0];
  assign mem_167_2_W0_clk = W0_clk;
  assign mem_167_2_W0_data = W0_data[23:16];
  assign mem_167_2_W0_en = W0_en & W0_addr_sel == 8'ha7;
  assign mem_167_2_W0_mask = W0_mask[2];
  assign mem_167_3_R0_addr = R0_addr[25:0];
  assign mem_167_3_R0_clk = R0_clk;
  assign mem_167_3_R0_en = R0_en & R0_addr_sel == 8'ha7;
  assign mem_167_3_W0_addr = W0_addr[25:0];
  assign mem_167_3_W0_clk = W0_clk;
  assign mem_167_3_W0_data = W0_data[31:24];
  assign mem_167_3_W0_en = W0_en & W0_addr_sel == 8'ha7;
  assign mem_167_3_W0_mask = W0_mask[3];
  assign mem_167_4_R0_addr = R0_addr[25:0];
  assign mem_167_4_R0_clk = R0_clk;
  assign mem_167_4_R0_en = R0_en & R0_addr_sel == 8'ha7;
  assign mem_167_4_W0_addr = W0_addr[25:0];
  assign mem_167_4_W0_clk = W0_clk;
  assign mem_167_4_W0_data = W0_data[39:32];
  assign mem_167_4_W0_en = W0_en & W0_addr_sel == 8'ha7;
  assign mem_167_4_W0_mask = W0_mask[4];
  assign mem_167_5_R0_addr = R0_addr[25:0];
  assign mem_167_5_R0_clk = R0_clk;
  assign mem_167_5_R0_en = R0_en & R0_addr_sel == 8'ha7;
  assign mem_167_5_W0_addr = W0_addr[25:0];
  assign mem_167_5_W0_clk = W0_clk;
  assign mem_167_5_W0_data = W0_data[47:40];
  assign mem_167_5_W0_en = W0_en & W0_addr_sel == 8'ha7;
  assign mem_167_5_W0_mask = W0_mask[5];
  assign mem_167_6_R0_addr = R0_addr[25:0];
  assign mem_167_6_R0_clk = R0_clk;
  assign mem_167_6_R0_en = R0_en & R0_addr_sel == 8'ha7;
  assign mem_167_6_W0_addr = W0_addr[25:0];
  assign mem_167_6_W0_clk = W0_clk;
  assign mem_167_6_W0_data = W0_data[55:48];
  assign mem_167_6_W0_en = W0_en & W0_addr_sel == 8'ha7;
  assign mem_167_6_W0_mask = W0_mask[6];
  assign mem_167_7_R0_addr = R0_addr[25:0];
  assign mem_167_7_R0_clk = R0_clk;
  assign mem_167_7_R0_en = R0_en & R0_addr_sel == 8'ha7;
  assign mem_167_7_W0_addr = W0_addr[25:0];
  assign mem_167_7_W0_clk = W0_clk;
  assign mem_167_7_W0_data = W0_data[63:56];
  assign mem_167_7_W0_en = W0_en & W0_addr_sel == 8'ha7;
  assign mem_167_7_W0_mask = W0_mask[7];
  assign mem_168_0_R0_addr = R0_addr[25:0];
  assign mem_168_0_R0_clk = R0_clk;
  assign mem_168_0_R0_en = R0_en & R0_addr_sel == 8'ha8;
  assign mem_168_0_W0_addr = W0_addr[25:0];
  assign mem_168_0_W0_clk = W0_clk;
  assign mem_168_0_W0_data = W0_data[7:0];
  assign mem_168_0_W0_en = W0_en & W0_addr_sel == 8'ha8;
  assign mem_168_0_W0_mask = W0_mask[0];
  assign mem_168_1_R0_addr = R0_addr[25:0];
  assign mem_168_1_R0_clk = R0_clk;
  assign mem_168_1_R0_en = R0_en & R0_addr_sel == 8'ha8;
  assign mem_168_1_W0_addr = W0_addr[25:0];
  assign mem_168_1_W0_clk = W0_clk;
  assign mem_168_1_W0_data = W0_data[15:8];
  assign mem_168_1_W0_en = W0_en & W0_addr_sel == 8'ha8;
  assign mem_168_1_W0_mask = W0_mask[1];
  assign mem_168_2_R0_addr = R0_addr[25:0];
  assign mem_168_2_R0_clk = R0_clk;
  assign mem_168_2_R0_en = R0_en & R0_addr_sel == 8'ha8;
  assign mem_168_2_W0_addr = W0_addr[25:0];
  assign mem_168_2_W0_clk = W0_clk;
  assign mem_168_2_W0_data = W0_data[23:16];
  assign mem_168_2_W0_en = W0_en & W0_addr_sel == 8'ha8;
  assign mem_168_2_W0_mask = W0_mask[2];
  assign mem_168_3_R0_addr = R0_addr[25:0];
  assign mem_168_3_R0_clk = R0_clk;
  assign mem_168_3_R0_en = R0_en & R0_addr_sel == 8'ha8;
  assign mem_168_3_W0_addr = W0_addr[25:0];
  assign mem_168_3_W0_clk = W0_clk;
  assign mem_168_3_W0_data = W0_data[31:24];
  assign mem_168_3_W0_en = W0_en & W0_addr_sel == 8'ha8;
  assign mem_168_3_W0_mask = W0_mask[3];
  assign mem_168_4_R0_addr = R0_addr[25:0];
  assign mem_168_4_R0_clk = R0_clk;
  assign mem_168_4_R0_en = R0_en & R0_addr_sel == 8'ha8;
  assign mem_168_4_W0_addr = W0_addr[25:0];
  assign mem_168_4_W0_clk = W0_clk;
  assign mem_168_4_W0_data = W0_data[39:32];
  assign mem_168_4_W0_en = W0_en & W0_addr_sel == 8'ha8;
  assign mem_168_4_W0_mask = W0_mask[4];
  assign mem_168_5_R0_addr = R0_addr[25:0];
  assign mem_168_5_R0_clk = R0_clk;
  assign mem_168_5_R0_en = R0_en & R0_addr_sel == 8'ha8;
  assign mem_168_5_W0_addr = W0_addr[25:0];
  assign mem_168_5_W0_clk = W0_clk;
  assign mem_168_5_W0_data = W0_data[47:40];
  assign mem_168_5_W0_en = W0_en & W0_addr_sel == 8'ha8;
  assign mem_168_5_W0_mask = W0_mask[5];
  assign mem_168_6_R0_addr = R0_addr[25:0];
  assign mem_168_6_R0_clk = R0_clk;
  assign mem_168_6_R0_en = R0_en & R0_addr_sel == 8'ha8;
  assign mem_168_6_W0_addr = W0_addr[25:0];
  assign mem_168_6_W0_clk = W0_clk;
  assign mem_168_6_W0_data = W0_data[55:48];
  assign mem_168_6_W0_en = W0_en & W0_addr_sel == 8'ha8;
  assign mem_168_6_W0_mask = W0_mask[6];
  assign mem_168_7_R0_addr = R0_addr[25:0];
  assign mem_168_7_R0_clk = R0_clk;
  assign mem_168_7_R0_en = R0_en & R0_addr_sel == 8'ha8;
  assign mem_168_7_W0_addr = W0_addr[25:0];
  assign mem_168_7_W0_clk = W0_clk;
  assign mem_168_7_W0_data = W0_data[63:56];
  assign mem_168_7_W0_en = W0_en & W0_addr_sel == 8'ha8;
  assign mem_168_7_W0_mask = W0_mask[7];
  assign mem_169_0_R0_addr = R0_addr[25:0];
  assign mem_169_0_R0_clk = R0_clk;
  assign mem_169_0_R0_en = R0_en & R0_addr_sel == 8'ha9;
  assign mem_169_0_W0_addr = W0_addr[25:0];
  assign mem_169_0_W0_clk = W0_clk;
  assign mem_169_0_W0_data = W0_data[7:0];
  assign mem_169_0_W0_en = W0_en & W0_addr_sel == 8'ha9;
  assign mem_169_0_W0_mask = W0_mask[0];
  assign mem_169_1_R0_addr = R0_addr[25:0];
  assign mem_169_1_R0_clk = R0_clk;
  assign mem_169_1_R0_en = R0_en & R0_addr_sel == 8'ha9;
  assign mem_169_1_W0_addr = W0_addr[25:0];
  assign mem_169_1_W0_clk = W0_clk;
  assign mem_169_1_W0_data = W0_data[15:8];
  assign mem_169_1_W0_en = W0_en & W0_addr_sel == 8'ha9;
  assign mem_169_1_W0_mask = W0_mask[1];
  assign mem_169_2_R0_addr = R0_addr[25:0];
  assign mem_169_2_R0_clk = R0_clk;
  assign mem_169_2_R0_en = R0_en & R0_addr_sel == 8'ha9;
  assign mem_169_2_W0_addr = W0_addr[25:0];
  assign mem_169_2_W0_clk = W0_clk;
  assign mem_169_2_W0_data = W0_data[23:16];
  assign mem_169_2_W0_en = W0_en & W0_addr_sel == 8'ha9;
  assign mem_169_2_W0_mask = W0_mask[2];
  assign mem_169_3_R0_addr = R0_addr[25:0];
  assign mem_169_3_R0_clk = R0_clk;
  assign mem_169_3_R0_en = R0_en & R0_addr_sel == 8'ha9;
  assign mem_169_3_W0_addr = W0_addr[25:0];
  assign mem_169_3_W0_clk = W0_clk;
  assign mem_169_3_W0_data = W0_data[31:24];
  assign mem_169_3_W0_en = W0_en & W0_addr_sel == 8'ha9;
  assign mem_169_3_W0_mask = W0_mask[3];
  assign mem_169_4_R0_addr = R0_addr[25:0];
  assign mem_169_4_R0_clk = R0_clk;
  assign mem_169_4_R0_en = R0_en & R0_addr_sel == 8'ha9;
  assign mem_169_4_W0_addr = W0_addr[25:0];
  assign mem_169_4_W0_clk = W0_clk;
  assign mem_169_4_W0_data = W0_data[39:32];
  assign mem_169_4_W0_en = W0_en & W0_addr_sel == 8'ha9;
  assign mem_169_4_W0_mask = W0_mask[4];
  assign mem_169_5_R0_addr = R0_addr[25:0];
  assign mem_169_5_R0_clk = R0_clk;
  assign mem_169_5_R0_en = R0_en & R0_addr_sel == 8'ha9;
  assign mem_169_5_W0_addr = W0_addr[25:0];
  assign mem_169_5_W0_clk = W0_clk;
  assign mem_169_5_W0_data = W0_data[47:40];
  assign mem_169_5_W0_en = W0_en & W0_addr_sel == 8'ha9;
  assign mem_169_5_W0_mask = W0_mask[5];
  assign mem_169_6_R0_addr = R0_addr[25:0];
  assign mem_169_6_R0_clk = R0_clk;
  assign mem_169_6_R0_en = R0_en & R0_addr_sel == 8'ha9;
  assign mem_169_6_W0_addr = W0_addr[25:0];
  assign mem_169_6_W0_clk = W0_clk;
  assign mem_169_6_W0_data = W0_data[55:48];
  assign mem_169_6_W0_en = W0_en & W0_addr_sel == 8'ha9;
  assign mem_169_6_W0_mask = W0_mask[6];
  assign mem_169_7_R0_addr = R0_addr[25:0];
  assign mem_169_7_R0_clk = R0_clk;
  assign mem_169_7_R0_en = R0_en & R0_addr_sel == 8'ha9;
  assign mem_169_7_W0_addr = W0_addr[25:0];
  assign mem_169_7_W0_clk = W0_clk;
  assign mem_169_7_W0_data = W0_data[63:56];
  assign mem_169_7_W0_en = W0_en & W0_addr_sel == 8'ha9;
  assign mem_169_7_W0_mask = W0_mask[7];
  assign mem_170_0_R0_addr = R0_addr[25:0];
  assign mem_170_0_R0_clk = R0_clk;
  assign mem_170_0_R0_en = R0_en & R0_addr_sel == 8'haa;
  assign mem_170_0_W0_addr = W0_addr[25:0];
  assign mem_170_0_W0_clk = W0_clk;
  assign mem_170_0_W0_data = W0_data[7:0];
  assign mem_170_0_W0_en = W0_en & W0_addr_sel == 8'haa;
  assign mem_170_0_W0_mask = W0_mask[0];
  assign mem_170_1_R0_addr = R0_addr[25:0];
  assign mem_170_1_R0_clk = R0_clk;
  assign mem_170_1_R0_en = R0_en & R0_addr_sel == 8'haa;
  assign mem_170_1_W0_addr = W0_addr[25:0];
  assign mem_170_1_W0_clk = W0_clk;
  assign mem_170_1_W0_data = W0_data[15:8];
  assign mem_170_1_W0_en = W0_en & W0_addr_sel == 8'haa;
  assign mem_170_1_W0_mask = W0_mask[1];
  assign mem_170_2_R0_addr = R0_addr[25:0];
  assign mem_170_2_R0_clk = R0_clk;
  assign mem_170_2_R0_en = R0_en & R0_addr_sel == 8'haa;
  assign mem_170_2_W0_addr = W0_addr[25:0];
  assign mem_170_2_W0_clk = W0_clk;
  assign mem_170_2_W0_data = W0_data[23:16];
  assign mem_170_2_W0_en = W0_en & W0_addr_sel == 8'haa;
  assign mem_170_2_W0_mask = W0_mask[2];
  assign mem_170_3_R0_addr = R0_addr[25:0];
  assign mem_170_3_R0_clk = R0_clk;
  assign mem_170_3_R0_en = R0_en & R0_addr_sel == 8'haa;
  assign mem_170_3_W0_addr = W0_addr[25:0];
  assign mem_170_3_W0_clk = W0_clk;
  assign mem_170_3_W0_data = W0_data[31:24];
  assign mem_170_3_W0_en = W0_en & W0_addr_sel == 8'haa;
  assign mem_170_3_W0_mask = W0_mask[3];
  assign mem_170_4_R0_addr = R0_addr[25:0];
  assign mem_170_4_R0_clk = R0_clk;
  assign mem_170_4_R0_en = R0_en & R0_addr_sel == 8'haa;
  assign mem_170_4_W0_addr = W0_addr[25:0];
  assign mem_170_4_W0_clk = W0_clk;
  assign mem_170_4_W0_data = W0_data[39:32];
  assign mem_170_4_W0_en = W0_en & W0_addr_sel == 8'haa;
  assign mem_170_4_W0_mask = W0_mask[4];
  assign mem_170_5_R0_addr = R0_addr[25:0];
  assign mem_170_5_R0_clk = R0_clk;
  assign mem_170_5_R0_en = R0_en & R0_addr_sel == 8'haa;
  assign mem_170_5_W0_addr = W0_addr[25:0];
  assign mem_170_5_W0_clk = W0_clk;
  assign mem_170_5_W0_data = W0_data[47:40];
  assign mem_170_5_W0_en = W0_en & W0_addr_sel == 8'haa;
  assign mem_170_5_W0_mask = W0_mask[5];
  assign mem_170_6_R0_addr = R0_addr[25:0];
  assign mem_170_6_R0_clk = R0_clk;
  assign mem_170_6_R0_en = R0_en & R0_addr_sel == 8'haa;
  assign mem_170_6_W0_addr = W0_addr[25:0];
  assign mem_170_6_W0_clk = W0_clk;
  assign mem_170_6_W0_data = W0_data[55:48];
  assign mem_170_6_W0_en = W0_en & W0_addr_sel == 8'haa;
  assign mem_170_6_W0_mask = W0_mask[6];
  assign mem_170_7_R0_addr = R0_addr[25:0];
  assign mem_170_7_R0_clk = R0_clk;
  assign mem_170_7_R0_en = R0_en & R0_addr_sel == 8'haa;
  assign mem_170_7_W0_addr = W0_addr[25:0];
  assign mem_170_7_W0_clk = W0_clk;
  assign mem_170_7_W0_data = W0_data[63:56];
  assign mem_170_7_W0_en = W0_en & W0_addr_sel == 8'haa;
  assign mem_170_7_W0_mask = W0_mask[7];
  assign mem_171_0_R0_addr = R0_addr[25:0];
  assign mem_171_0_R0_clk = R0_clk;
  assign mem_171_0_R0_en = R0_en & R0_addr_sel == 8'hab;
  assign mem_171_0_W0_addr = W0_addr[25:0];
  assign mem_171_0_W0_clk = W0_clk;
  assign mem_171_0_W0_data = W0_data[7:0];
  assign mem_171_0_W0_en = W0_en & W0_addr_sel == 8'hab;
  assign mem_171_0_W0_mask = W0_mask[0];
  assign mem_171_1_R0_addr = R0_addr[25:0];
  assign mem_171_1_R0_clk = R0_clk;
  assign mem_171_1_R0_en = R0_en & R0_addr_sel == 8'hab;
  assign mem_171_1_W0_addr = W0_addr[25:0];
  assign mem_171_1_W0_clk = W0_clk;
  assign mem_171_1_W0_data = W0_data[15:8];
  assign mem_171_1_W0_en = W0_en & W0_addr_sel == 8'hab;
  assign mem_171_1_W0_mask = W0_mask[1];
  assign mem_171_2_R0_addr = R0_addr[25:0];
  assign mem_171_2_R0_clk = R0_clk;
  assign mem_171_2_R0_en = R0_en & R0_addr_sel == 8'hab;
  assign mem_171_2_W0_addr = W0_addr[25:0];
  assign mem_171_2_W0_clk = W0_clk;
  assign mem_171_2_W0_data = W0_data[23:16];
  assign mem_171_2_W0_en = W0_en & W0_addr_sel == 8'hab;
  assign mem_171_2_W0_mask = W0_mask[2];
  assign mem_171_3_R0_addr = R0_addr[25:0];
  assign mem_171_3_R0_clk = R0_clk;
  assign mem_171_3_R0_en = R0_en & R0_addr_sel == 8'hab;
  assign mem_171_3_W0_addr = W0_addr[25:0];
  assign mem_171_3_W0_clk = W0_clk;
  assign mem_171_3_W0_data = W0_data[31:24];
  assign mem_171_3_W0_en = W0_en & W0_addr_sel == 8'hab;
  assign mem_171_3_W0_mask = W0_mask[3];
  assign mem_171_4_R0_addr = R0_addr[25:0];
  assign mem_171_4_R0_clk = R0_clk;
  assign mem_171_4_R0_en = R0_en & R0_addr_sel == 8'hab;
  assign mem_171_4_W0_addr = W0_addr[25:0];
  assign mem_171_4_W0_clk = W0_clk;
  assign mem_171_4_W0_data = W0_data[39:32];
  assign mem_171_4_W0_en = W0_en & W0_addr_sel == 8'hab;
  assign mem_171_4_W0_mask = W0_mask[4];
  assign mem_171_5_R0_addr = R0_addr[25:0];
  assign mem_171_5_R0_clk = R0_clk;
  assign mem_171_5_R0_en = R0_en & R0_addr_sel == 8'hab;
  assign mem_171_5_W0_addr = W0_addr[25:0];
  assign mem_171_5_W0_clk = W0_clk;
  assign mem_171_5_W0_data = W0_data[47:40];
  assign mem_171_5_W0_en = W0_en & W0_addr_sel == 8'hab;
  assign mem_171_5_W0_mask = W0_mask[5];
  assign mem_171_6_R0_addr = R0_addr[25:0];
  assign mem_171_6_R0_clk = R0_clk;
  assign mem_171_6_R0_en = R0_en & R0_addr_sel == 8'hab;
  assign mem_171_6_W0_addr = W0_addr[25:0];
  assign mem_171_6_W0_clk = W0_clk;
  assign mem_171_6_W0_data = W0_data[55:48];
  assign mem_171_6_W0_en = W0_en & W0_addr_sel == 8'hab;
  assign mem_171_6_W0_mask = W0_mask[6];
  assign mem_171_7_R0_addr = R0_addr[25:0];
  assign mem_171_7_R0_clk = R0_clk;
  assign mem_171_7_R0_en = R0_en & R0_addr_sel == 8'hab;
  assign mem_171_7_W0_addr = W0_addr[25:0];
  assign mem_171_7_W0_clk = W0_clk;
  assign mem_171_7_W0_data = W0_data[63:56];
  assign mem_171_7_W0_en = W0_en & W0_addr_sel == 8'hab;
  assign mem_171_7_W0_mask = W0_mask[7];
  assign mem_172_0_R0_addr = R0_addr[25:0];
  assign mem_172_0_R0_clk = R0_clk;
  assign mem_172_0_R0_en = R0_en & R0_addr_sel == 8'hac;
  assign mem_172_0_W0_addr = W0_addr[25:0];
  assign mem_172_0_W0_clk = W0_clk;
  assign mem_172_0_W0_data = W0_data[7:0];
  assign mem_172_0_W0_en = W0_en & W0_addr_sel == 8'hac;
  assign mem_172_0_W0_mask = W0_mask[0];
  assign mem_172_1_R0_addr = R0_addr[25:0];
  assign mem_172_1_R0_clk = R0_clk;
  assign mem_172_1_R0_en = R0_en & R0_addr_sel == 8'hac;
  assign mem_172_1_W0_addr = W0_addr[25:0];
  assign mem_172_1_W0_clk = W0_clk;
  assign mem_172_1_W0_data = W0_data[15:8];
  assign mem_172_1_W0_en = W0_en & W0_addr_sel == 8'hac;
  assign mem_172_1_W0_mask = W0_mask[1];
  assign mem_172_2_R0_addr = R0_addr[25:0];
  assign mem_172_2_R0_clk = R0_clk;
  assign mem_172_2_R0_en = R0_en & R0_addr_sel == 8'hac;
  assign mem_172_2_W0_addr = W0_addr[25:0];
  assign mem_172_2_W0_clk = W0_clk;
  assign mem_172_2_W0_data = W0_data[23:16];
  assign mem_172_2_W0_en = W0_en & W0_addr_sel == 8'hac;
  assign mem_172_2_W0_mask = W0_mask[2];
  assign mem_172_3_R0_addr = R0_addr[25:0];
  assign mem_172_3_R0_clk = R0_clk;
  assign mem_172_3_R0_en = R0_en & R0_addr_sel == 8'hac;
  assign mem_172_3_W0_addr = W0_addr[25:0];
  assign mem_172_3_W0_clk = W0_clk;
  assign mem_172_3_W0_data = W0_data[31:24];
  assign mem_172_3_W0_en = W0_en & W0_addr_sel == 8'hac;
  assign mem_172_3_W0_mask = W0_mask[3];
  assign mem_172_4_R0_addr = R0_addr[25:0];
  assign mem_172_4_R0_clk = R0_clk;
  assign mem_172_4_R0_en = R0_en & R0_addr_sel == 8'hac;
  assign mem_172_4_W0_addr = W0_addr[25:0];
  assign mem_172_4_W0_clk = W0_clk;
  assign mem_172_4_W0_data = W0_data[39:32];
  assign mem_172_4_W0_en = W0_en & W0_addr_sel == 8'hac;
  assign mem_172_4_W0_mask = W0_mask[4];
  assign mem_172_5_R0_addr = R0_addr[25:0];
  assign mem_172_5_R0_clk = R0_clk;
  assign mem_172_5_R0_en = R0_en & R0_addr_sel == 8'hac;
  assign mem_172_5_W0_addr = W0_addr[25:0];
  assign mem_172_5_W0_clk = W0_clk;
  assign mem_172_5_W0_data = W0_data[47:40];
  assign mem_172_5_W0_en = W0_en & W0_addr_sel == 8'hac;
  assign mem_172_5_W0_mask = W0_mask[5];
  assign mem_172_6_R0_addr = R0_addr[25:0];
  assign mem_172_6_R0_clk = R0_clk;
  assign mem_172_6_R0_en = R0_en & R0_addr_sel == 8'hac;
  assign mem_172_6_W0_addr = W0_addr[25:0];
  assign mem_172_6_W0_clk = W0_clk;
  assign mem_172_6_W0_data = W0_data[55:48];
  assign mem_172_6_W0_en = W0_en & W0_addr_sel == 8'hac;
  assign mem_172_6_W0_mask = W0_mask[6];
  assign mem_172_7_R0_addr = R0_addr[25:0];
  assign mem_172_7_R0_clk = R0_clk;
  assign mem_172_7_R0_en = R0_en & R0_addr_sel == 8'hac;
  assign mem_172_7_W0_addr = W0_addr[25:0];
  assign mem_172_7_W0_clk = W0_clk;
  assign mem_172_7_W0_data = W0_data[63:56];
  assign mem_172_7_W0_en = W0_en & W0_addr_sel == 8'hac;
  assign mem_172_7_W0_mask = W0_mask[7];
  assign mem_173_0_R0_addr = R0_addr[25:0];
  assign mem_173_0_R0_clk = R0_clk;
  assign mem_173_0_R0_en = R0_en & R0_addr_sel == 8'had;
  assign mem_173_0_W0_addr = W0_addr[25:0];
  assign mem_173_0_W0_clk = W0_clk;
  assign mem_173_0_W0_data = W0_data[7:0];
  assign mem_173_0_W0_en = W0_en & W0_addr_sel == 8'had;
  assign mem_173_0_W0_mask = W0_mask[0];
  assign mem_173_1_R0_addr = R0_addr[25:0];
  assign mem_173_1_R0_clk = R0_clk;
  assign mem_173_1_R0_en = R0_en & R0_addr_sel == 8'had;
  assign mem_173_1_W0_addr = W0_addr[25:0];
  assign mem_173_1_W0_clk = W0_clk;
  assign mem_173_1_W0_data = W0_data[15:8];
  assign mem_173_1_W0_en = W0_en & W0_addr_sel == 8'had;
  assign mem_173_1_W0_mask = W0_mask[1];
  assign mem_173_2_R0_addr = R0_addr[25:0];
  assign mem_173_2_R0_clk = R0_clk;
  assign mem_173_2_R0_en = R0_en & R0_addr_sel == 8'had;
  assign mem_173_2_W0_addr = W0_addr[25:0];
  assign mem_173_2_W0_clk = W0_clk;
  assign mem_173_2_W0_data = W0_data[23:16];
  assign mem_173_2_W0_en = W0_en & W0_addr_sel == 8'had;
  assign mem_173_2_W0_mask = W0_mask[2];
  assign mem_173_3_R0_addr = R0_addr[25:0];
  assign mem_173_3_R0_clk = R0_clk;
  assign mem_173_3_R0_en = R0_en & R0_addr_sel == 8'had;
  assign mem_173_3_W0_addr = W0_addr[25:0];
  assign mem_173_3_W0_clk = W0_clk;
  assign mem_173_3_W0_data = W0_data[31:24];
  assign mem_173_3_W0_en = W0_en & W0_addr_sel == 8'had;
  assign mem_173_3_W0_mask = W0_mask[3];
  assign mem_173_4_R0_addr = R0_addr[25:0];
  assign mem_173_4_R0_clk = R0_clk;
  assign mem_173_4_R0_en = R0_en & R0_addr_sel == 8'had;
  assign mem_173_4_W0_addr = W0_addr[25:0];
  assign mem_173_4_W0_clk = W0_clk;
  assign mem_173_4_W0_data = W0_data[39:32];
  assign mem_173_4_W0_en = W0_en & W0_addr_sel == 8'had;
  assign mem_173_4_W0_mask = W0_mask[4];
  assign mem_173_5_R0_addr = R0_addr[25:0];
  assign mem_173_5_R0_clk = R0_clk;
  assign mem_173_5_R0_en = R0_en & R0_addr_sel == 8'had;
  assign mem_173_5_W0_addr = W0_addr[25:0];
  assign mem_173_5_W0_clk = W0_clk;
  assign mem_173_5_W0_data = W0_data[47:40];
  assign mem_173_5_W0_en = W0_en & W0_addr_sel == 8'had;
  assign mem_173_5_W0_mask = W0_mask[5];
  assign mem_173_6_R0_addr = R0_addr[25:0];
  assign mem_173_6_R0_clk = R0_clk;
  assign mem_173_6_R0_en = R0_en & R0_addr_sel == 8'had;
  assign mem_173_6_W0_addr = W0_addr[25:0];
  assign mem_173_6_W0_clk = W0_clk;
  assign mem_173_6_W0_data = W0_data[55:48];
  assign mem_173_6_W0_en = W0_en & W0_addr_sel == 8'had;
  assign mem_173_6_W0_mask = W0_mask[6];
  assign mem_173_7_R0_addr = R0_addr[25:0];
  assign mem_173_7_R0_clk = R0_clk;
  assign mem_173_7_R0_en = R0_en & R0_addr_sel == 8'had;
  assign mem_173_7_W0_addr = W0_addr[25:0];
  assign mem_173_7_W0_clk = W0_clk;
  assign mem_173_7_W0_data = W0_data[63:56];
  assign mem_173_7_W0_en = W0_en & W0_addr_sel == 8'had;
  assign mem_173_7_W0_mask = W0_mask[7];
  assign mem_174_0_R0_addr = R0_addr[25:0];
  assign mem_174_0_R0_clk = R0_clk;
  assign mem_174_0_R0_en = R0_en & R0_addr_sel == 8'hae;
  assign mem_174_0_W0_addr = W0_addr[25:0];
  assign mem_174_0_W0_clk = W0_clk;
  assign mem_174_0_W0_data = W0_data[7:0];
  assign mem_174_0_W0_en = W0_en & W0_addr_sel == 8'hae;
  assign mem_174_0_W0_mask = W0_mask[0];
  assign mem_174_1_R0_addr = R0_addr[25:0];
  assign mem_174_1_R0_clk = R0_clk;
  assign mem_174_1_R0_en = R0_en & R0_addr_sel == 8'hae;
  assign mem_174_1_W0_addr = W0_addr[25:0];
  assign mem_174_1_W0_clk = W0_clk;
  assign mem_174_1_W0_data = W0_data[15:8];
  assign mem_174_1_W0_en = W0_en & W0_addr_sel == 8'hae;
  assign mem_174_1_W0_mask = W0_mask[1];
  assign mem_174_2_R0_addr = R0_addr[25:0];
  assign mem_174_2_R0_clk = R0_clk;
  assign mem_174_2_R0_en = R0_en & R0_addr_sel == 8'hae;
  assign mem_174_2_W0_addr = W0_addr[25:0];
  assign mem_174_2_W0_clk = W0_clk;
  assign mem_174_2_W0_data = W0_data[23:16];
  assign mem_174_2_W0_en = W0_en & W0_addr_sel == 8'hae;
  assign mem_174_2_W0_mask = W0_mask[2];
  assign mem_174_3_R0_addr = R0_addr[25:0];
  assign mem_174_3_R0_clk = R0_clk;
  assign mem_174_3_R0_en = R0_en & R0_addr_sel == 8'hae;
  assign mem_174_3_W0_addr = W0_addr[25:0];
  assign mem_174_3_W0_clk = W0_clk;
  assign mem_174_3_W0_data = W0_data[31:24];
  assign mem_174_3_W0_en = W0_en & W0_addr_sel == 8'hae;
  assign mem_174_3_W0_mask = W0_mask[3];
  assign mem_174_4_R0_addr = R0_addr[25:0];
  assign mem_174_4_R0_clk = R0_clk;
  assign mem_174_4_R0_en = R0_en & R0_addr_sel == 8'hae;
  assign mem_174_4_W0_addr = W0_addr[25:0];
  assign mem_174_4_W0_clk = W0_clk;
  assign mem_174_4_W0_data = W0_data[39:32];
  assign mem_174_4_W0_en = W0_en & W0_addr_sel == 8'hae;
  assign mem_174_4_W0_mask = W0_mask[4];
  assign mem_174_5_R0_addr = R0_addr[25:0];
  assign mem_174_5_R0_clk = R0_clk;
  assign mem_174_5_R0_en = R0_en & R0_addr_sel == 8'hae;
  assign mem_174_5_W0_addr = W0_addr[25:0];
  assign mem_174_5_W0_clk = W0_clk;
  assign mem_174_5_W0_data = W0_data[47:40];
  assign mem_174_5_W0_en = W0_en & W0_addr_sel == 8'hae;
  assign mem_174_5_W0_mask = W0_mask[5];
  assign mem_174_6_R0_addr = R0_addr[25:0];
  assign mem_174_6_R0_clk = R0_clk;
  assign mem_174_6_R0_en = R0_en & R0_addr_sel == 8'hae;
  assign mem_174_6_W0_addr = W0_addr[25:0];
  assign mem_174_6_W0_clk = W0_clk;
  assign mem_174_6_W0_data = W0_data[55:48];
  assign mem_174_6_W0_en = W0_en & W0_addr_sel == 8'hae;
  assign mem_174_6_W0_mask = W0_mask[6];
  assign mem_174_7_R0_addr = R0_addr[25:0];
  assign mem_174_7_R0_clk = R0_clk;
  assign mem_174_7_R0_en = R0_en & R0_addr_sel == 8'hae;
  assign mem_174_7_W0_addr = W0_addr[25:0];
  assign mem_174_7_W0_clk = W0_clk;
  assign mem_174_7_W0_data = W0_data[63:56];
  assign mem_174_7_W0_en = W0_en & W0_addr_sel == 8'hae;
  assign mem_174_7_W0_mask = W0_mask[7];
  assign mem_175_0_R0_addr = R0_addr[25:0];
  assign mem_175_0_R0_clk = R0_clk;
  assign mem_175_0_R0_en = R0_en & R0_addr_sel == 8'haf;
  assign mem_175_0_W0_addr = W0_addr[25:0];
  assign mem_175_0_W0_clk = W0_clk;
  assign mem_175_0_W0_data = W0_data[7:0];
  assign mem_175_0_W0_en = W0_en & W0_addr_sel == 8'haf;
  assign mem_175_0_W0_mask = W0_mask[0];
  assign mem_175_1_R0_addr = R0_addr[25:0];
  assign mem_175_1_R0_clk = R0_clk;
  assign mem_175_1_R0_en = R0_en & R0_addr_sel == 8'haf;
  assign mem_175_1_W0_addr = W0_addr[25:0];
  assign mem_175_1_W0_clk = W0_clk;
  assign mem_175_1_W0_data = W0_data[15:8];
  assign mem_175_1_W0_en = W0_en & W0_addr_sel == 8'haf;
  assign mem_175_1_W0_mask = W0_mask[1];
  assign mem_175_2_R0_addr = R0_addr[25:0];
  assign mem_175_2_R0_clk = R0_clk;
  assign mem_175_2_R0_en = R0_en & R0_addr_sel == 8'haf;
  assign mem_175_2_W0_addr = W0_addr[25:0];
  assign mem_175_2_W0_clk = W0_clk;
  assign mem_175_2_W0_data = W0_data[23:16];
  assign mem_175_2_W0_en = W0_en & W0_addr_sel == 8'haf;
  assign mem_175_2_W0_mask = W0_mask[2];
  assign mem_175_3_R0_addr = R0_addr[25:0];
  assign mem_175_3_R0_clk = R0_clk;
  assign mem_175_3_R0_en = R0_en & R0_addr_sel == 8'haf;
  assign mem_175_3_W0_addr = W0_addr[25:0];
  assign mem_175_3_W0_clk = W0_clk;
  assign mem_175_3_W0_data = W0_data[31:24];
  assign mem_175_3_W0_en = W0_en & W0_addr_sel == 8'haf;
  assign mem_175_3_W0_mask = W0_mask[3];
  assign mem_175_4_R0_addr = R0_addr[25:0];
  assign mem_175_4_R0_clk = R0_clk;
  assign mem_175_4_R0_en = R0_en & R0_addr_sel == 8'haf;
  assign mem_175_4_W0_addr = W0_addr[25:0];
  assign mem_175_4_W0_clk = W0_clk;
  assign mem_175_4_W0_data = W0_data[39:32];
  assign mem_175_4_W0_en = W0_en & W0_addr_sel == 8'haf;
  assign mem_175_4_W0_mask = W0_mask[4];
  assign mem_175_5_R0_addr = R0_addr[25:0];
  assign mem_175_5_R0_clk = R0_clk;
  assign mem_175_5_R0_en = R0_en & R0_addr_sel == 8'haf;
  assign mem_175_5_W0_addr = W0_addr[25:0];
  assign mem_175_5_W0_clk = W0_clk;
  assign mem_175_5_W0_data = W0_data[47:40];
  assign mem_175_5_W0_en = W0_en & W0_addr_sel == 8'haf;
  assign mem_175_5_W0_mask = W0_mask[5];
  assign mem_175_6_R0_addr = R0_addr[25:0];
  assign mem_175_6_R0_clk = R0_clk;
  assign mem_175_6_R0_en = R0_en & R0_addr_sel == 8'haf;
  assign mem_175_6_W0_addr = W0_addr[25:0];
  assign mem_175_6_W0_clk = W0_clk;
  assign mem_175_6_W0_data = W0_data[55:48];
  assign mem_175_6_W0_en = W0_en & W0_addr_sel == 8'haf;
  assign mem_175_6_W0_mask = W0_mask[6];
  assign mem_175_7_R0_addr = R0_addr[25:0];
  assign mem_175_7_R0_clk = R0_clk;
  assign mem_175_7_R0_en = R0_en & R0_addr_sel == 8'haf;
  assign mem_175_7_W0_addr = W0_addr[25:0];
  assign mem_175_7_W0_clk = W0_clk;
  assign mem_175_7_W0_data = W0_data[63:56];
  assign mem_175_7_W0_en = W0_en & W0_addr_sel == 8'haf;
  assign mem_175_7_W0_mask = W0_mask[7];
  assign mem_176_0_R0_addr = R0_addr[25:0];
  assign mem_176_0_R0_clk = R0_clk;
  assign mem_176_0_R0_en = R0_en & R0_addr_sel == 8'hb0;
  assign mem_176_0_W0_addr = W0_addr[25:0];
  assign mem_176_0_W0_clk = W0_clk;
  assign mem_176_0_W0_data = W0_data[7:0];
  assign mem_176_0_W0_en = W0_en & W0_addr_sel == 8'hb0;
  assign mem_176_0_W0_mask = W0_mask[0];
  assign mem_176_1_R0_addr = R0_addr[25:0];
  assign mem_176_1_R0_clk = R0_clk;
  assign mem_176_1_R0_en = R0_en & R0_addr_sel == 8'hb0;
  assign mem_176_1_W0_addr = W0_addr[25:0];
  assign mem_176_1_W0_clk = W0_clk;
  assign mem_176_1_W0_data = W0_data[15:8];
  assign mem_176_1_W0_en = W0_en & W0_addr_sel == 8'hb0;
  assign mem_176_1_W0_mask = W0_mask[1];
  assign mem_176_2_R0_addr = R0_addr[25:0];
  assign mem_176_2_R0_clk = R0_clk;
  assign mem_176_2_R0_en = R0_en & R0_addr_sel == 8'hb0;
  assign mem_176_2_W0_addr = W0_addr[25:0];
  assign mem_176_2_W0_clk = W0_clk;
  assign mem_176_2_W0_data = W0_data[23:16];
  assign mem_176_2_W0_en = W0_en & W0_addr_sel == 8'hb0;
  assign mem_176_2_W0_mask = W0_mask[2];
  assign mem_176_3_R0_addr = R0_addr[25:0];
  assign mem_176_3_R0_clk = R0_clk;
  assign mem_176_3_R0_en = R0_en & R0_addr_sel == 8'hb0;
  assign mem_176_3_W0_addr = W0_addr[25:0];
  assign mem_176_3_W0_clk = W0_clk;
  assign mem_176_3_W0_data = W0_data[31:24];
  assign mem_176_3_W0_en = W0_en & W0_addr_sel == 8'hb0;
  assign mem_176_3_W0_mask = W0_mask[3];
  assign mem_176_4_R0_addr = R0_addr[25:0];
  assign mem_176_4_R0_clk = R0_clk;
  assign mem_176_4_R0_en = R0_en & R0_addr_sel == 8'hb0;
  assign mem_176_4_W0_addr = W0_addr[25:0];
  assign mem_176_4_W0_clk = W0_clk;
  assign mem_176_4_W0_data = W0_data[39:32];
  assign mem_176_4_W0_en = W0_en & W0_addr_sel == 8'hb0;
  assign mem_176_4_W0_mask = W0_mask[4];
  assign mem_176_5_R0_addr = R0_addr[25:0];
  assign mem_176_5_R0_clk = R0_clk;
  assign mem_176_5_R0_en = R0_en & R0_addr_sel == 8'hb0;
  assign mem_176_5_W0_addr = W0_addr[25:0];
  assign mem_176_5_W0_clk = W0_clk;
  assign mem_176_5_W0_data = W0_data[47:40];
  assign mem_176_5_W0_en = W0_en & W0_addr_sel == 8'hb0;
  assign mem_176_5_W0_mask = W0_mask[5];
  assign mem_176_6_R0_addr = R0_addr[25:0];
  assign mem_176_6_R0_clk = R0_clk;
  assign mem_176_6_R0_en = R0_en & R0_addr_sel == 8'hb0;
  assign mem_176_6_W0_addr = W0_addr[25:0];
  assign mem_176_6_W0_clk = W0_clk;
  assign mem_176_6_W0_data = W0_data[55:48];
  assign mem_176_6_W0_en = W0_en & W0_addr_sel == 8'hb0;
  assign mem_176_6_W0_mask = W0_mask[6];
  assign mem_176_7_R0_addr = R0_addr[25:0];
  assign mem_176_7_R0_clk = R0_clk;
  assign mem_176_7_R0_en = R0_en & R0_addr_sel == 8'hb0;
  assign mem_176_7_W0_addr = W0_addr[25:0];
  assign mem_176_7_W0_clk = W0_clk;
  assign mem_176_7_W0_data = W0_data[63:56];
  assign mem_176_7_W0_en = W0_en & W0_addr_sel == 8'hb0;
  assign mem_176_7_W0_mask = W0_mask[7];
  assign mem_177_0_R0_addr = R0_addr[25:0];
  assign mem_177_0_R0_clk = R0_clk;
  assign mem_177_0_R0_en = R0_en & R0_addr_sel == 8'hb1;
  assign mem_177_0_W0_addr = W0_addr[25:0];
  assign mem_177_0_W0_clk = W0_clk;
  assign mem_177_0_W0_data = W0_data[7:0];
  assign mem_177_0_W0_en = W0_en & W0_addr_sel == 8'hb1;
  assign mem_177_0_W0_mask = W0_mask[0];
  assign mem_177_1_R0_addr = R0_addr[25:0];
  assign mem_177_1_R0_clk = R0_clk;
  assign mem_177_1_R0_en = R0_en & R0_addr_sel == 8'hb1;
  assign mem_177_1_W0_addr = W0_addr[25:0];
  assign mem_177_1_W0_clk = W0_clk;
  assign mem_177_1_W0_data = W0_data[15:8];
  assign mem_177_1_W0_en = W0_en & W0_addr_sel == 8'hb1;
  assign mem_177_1_W0_mask = W0_mask[1];
  assign mem_177_2_R0_addr = R0_addr[25:0];
  assign mem_177_2_R0_clk = R0_clk;
  assign mem_177_2_R0_en = R0_en & R0_addr_sel == 8'hb1;
  assign mem_177_2_W0_addr = W0_addr[25:0];
  assign mem_177_2_W0_clk = W0_clk;
  assign mem_177_2_W0_data = W0_data[23:16];
  assign mem_177_2_W0_en = W0_en & W0_addr_sel == 8'hb1;
  assign mem_177_2_W0_mask = W0_mask[2];
  assign mem_177_3_R0_addr = R0_addr[25:0];
  assign mem_177_3_R0_clk = R0_clk;
  assign mem_177_3_R0_en = R0_en & R0_addr_sel == 8'hb1;
  assign mem_177_3_W0_addr = W0_addr[25:0];
  assign mem_177_3_W0_clk = W0_clk;
  assign mem_177_3_W0_data = W0_data[31:24];
  assign mem_177_3_W0_en = W0_en & W0_addr_sel == 8'hb1;
  assign mem_177_3_W0_mask = W0_mask[3];
  assign mem_177_4_R0_addr = R0_addr[25:0];
  assign mem_177_4_R0_clk = R0_clk;
  assign mem_177_4_R0_en = R0_en & R0_addr_sel == 8'hb1;
  assign mem_177_4_W0_addr = W0_addr[25:0];
  assign mem_177_4_W0_clk = W0_clk;
  assign mem_177_4_W0_data = W0_data[39:32];
  assign mem_177_4_W0_en = W0_en & W0_addr_sel == 8'hb1;
  assign mem_177_4_W0_mask = W0_mask[4];
  assign mem_177_5_R0_addr = R0_addr[25:0];
  assign mem_177_5_R0_clk = R0_clk;
  assign mem_177_5_R0_en = R0_en & R0_addr_sel == 8'hb1;
  assign mem_177_5_W0_addr = W0_addr[25:0];
  assign mem_177_5_W0_clk = W0_clk;
  assign mem_177_5_W0_data = W0_data[47:40];
  assign mem_177_5_W0_en = W0_en & W0_addr_sel == 8'hb1;
  assign mem_177_5_W0_mask = W0_mask[5];
  assign mem_177_6_R0_addr = R0_addr[25:0];
  assign mem_177_6_R0_clk = R0_clk;
  assign mem_177_6_R0_en = R0_en & R0_addr_sel == 8'hb1;
  assign mem_177_6_W0_addr = W0_addr[25:0];
  assign mem_177_6_W0_clk = W0_clk;
  assign mem_177_6_W0_data = W0_data[55:48];
  assign mem_177_6_W0_en = W0_en & W0_addr_sel == 8'hb1;
  assign mem_177_6_W0_mask = W0_mask[6];
  assign mem_177_7_R0_addr = R0_addr[25:0];
  assign mem_177_7_R0_clk = R0_clk;
  assign mem_177_7_R0_en = R0_en & R0_addr_sel == 8'hb1;
  assign mem_177_7_W0_addr = W0_addr[25:0];
  assign mem_177_7_W0_clk = W0_clk;
  assign mem_177_7_W0_data = W0_data[63:56];
  assign mem_177_7_W0_en = W0_en & W0_addr_sel == 8'hb1;
  assign mem_177_7_W0_mask = W0_mask[7];
  assign mem_178_0_R0_addr = R0_addr[25:0];
  assign mem_178_0_R0_clk = R0_clk;
  assign mem_178_0_R0_en = R0_en & R0_addr_sel == 8'hb2;
  assign mem_178_0_W0_addr = W0_addr[25:0];
  assign mem_178_0_W0_clk = W0_clk;
  assign mem_178_0_W0_data = W0_data[7:0];
  assign mem_178_0_W0_en = W0_en & W0_addr_sel == 8'hb2;
  assign mem_178_0_W0_mask = W0_mask[0];
  assign mem_178_1_R0_addr = R0_addr[25:0];
  assign mem_178_1_R0_clk = R0_clk;
  assign mem_178_1_R0_en = R0_en & R0_addr_sel == 8'hb2;
  assign mem_178_1_W0_addr = W0_addr[25:0];
  assign mem_178_1_W0_clk = W0_clk;
  assign mem_178_1_W0_data = W0_data[15:8];
  assign mem_178_1_W0_en = W0_en & W0_addr_sel == 8'hb2;
  assign mem_178_1_W0_mask = W0_mask[1];
  assign mem_178_2_R0_addr = R0_addr[25:0];
  assign mem_178_2_R0_clk = R0_clk;
  assign mem_178_2_R0_en = R0_en & R0_addr_sel == 8'hb2;
  assign mem_178_2_W0_addr = W0_addr[25:0];
  assign mem_178_2_W0_clk = W0_clk;
  assign mem_178_2_W0_data = W0_data[23:16];
  assign mem_178_2_W0_en = W0_en & W0_addr_sel == 8'hb2;
  assign mem_178_2_W0_mask = W0_mask[2];
  assign mem_178_3_R0_addr = R0_addr[25:0];
  assign mem_178_3_R0_clk = R0_clk;
  assign mem_178_3_R0_en = R0_en & R0_addr_sel == 8'hb2;
  assign mem_178_3_W0_addr = W0_addr[25:0];
  assign mem_178_3_W0_clk = W0_clk;
  assign mem_178_3_W0_data = W0_data[31:24];
  assign mem_178_3_W0_en = W0_en & W0_addr_sel == 8'hb2;
  assign mem_178_3_W0_mask = W0_mask[3];
  assign mem_178_4_R0_addr = R0_addr[25:0];
  assign mem_178_4_R0_clk = R0_clk;
  assign mem_178_4_R0_en = R0_en & R0_addr_sel == 8'hb2;
  assign mem_178_4_W0_addr = W0_addr[25:0];
  assign mem_178_4_W0_clk = W0_clk;
  assign mem_178_4_W0_data = W0_data[39:32];
  assign mem_178_4_W0_en = W0_en & W0_addr_sel == 8'hb2;
  assign mem_178_4_W0_mask = W0_mask[4];
  assign mem_178_5_R0_addr = R0_addr[25:0];
  assign mem_178_5_R0_clk = R0_clk;
  assign mem_178_5_R0_en = R0_en & R0_addr_sel == 8'hb2;
  assign mem_178_5_W0_addr = W0_addr[25:0];
  assign mem_178_5_W0_clk = W0_clk;
  assign mem_178_5_W0_data = W0_data[47:40];
  assign mem_178_5_W0_en = W0_en & W0_addr_sel == 8'hb2;
  assign mem_178_5_W0_mask = W0_mask[5];
  assign mem_178_6_R0_addr = R0_addr[25:0];
  assign mem_178_6_R0_clk = R0_clk;
  assign mem_178_6_R0_en = R0_en & R0_addr_sel == 8'hb2;
  assign mem_178_6_W0_addr = W0_addr[25:0];
  assign mem_178_6_W0_clk = W0_clk;
  assign mem_178_6_W0_data = W0_data[55:48];
  assign mem_178_6_W0_en = W0_en & W0_addr_sel == 8'hb2;
  assign mem_178_6_W0_mask = W0_mask[6];
  assign mem_178_7_R0_addr = R0_addr[25:0];
  assign mem_178_7_R0_clk = R0_clk;
  assign mem_178_7_R0_en = R0_en & R0_addr_sel == 8'hb2;
  assign mem_178_7_W0_addr = W0_addr[25:0];
  assign mem_178_7_W0_clk = W0_clk;
  assign mem_178_7_W0_data = W0_data[63:56];
  assign mem_178_7_W0_en = W0_en & W0_addr_sel == 8'hb2;
  assign mem_178_7_W0_mask = W0_mask[7];
  assign mem_179_0_R0_addr = R0_addr[25:0];
  assign mem_179_0_R0_clk = R0_clk;
  assign mem_179_0_R0_en = R0_en & R0_addr_sel == 8'hb3;
  assign mem_179_0_W0_addr = W0_addr[25:0];
  assign mem_179_0_W0_clk = W0_clk;
  assign mem_179_0_W0_data = W0_data[7:0];
  assign mem_179_0_W0_en = W0_en & W0_addr_sel == 8'hb3;
  assign mem_179_0_W0_mask = W0_mask[0];
  assign mem_179_1_R0_addr = R0_addr[25:0];
  assign mem_179_1_R0_clk = R0_clk;
  assign mem_179_1_R0_en = R0_en & R0_addr_sel == 8'hb3;
  assign mem_179_1_W0_addr = W0_addr[25:0];
  assign mem_179_1_W0_clk = W0_clk;
  assign mem_179_1_W0_data = W0_data[15:8];
  assign mem_179_1_W0_en = W0_en & W0_addr_sel == 8'hb3;
  assign mem_179_1_W0_mask = W0_mask[1];
  assign mem_179_2_R0_addr = R0_addr[25:0];
  assign mem_179_2_R0_clk = R0_clk;
  assign mem_179_2_R0_en = R0_en & R0_addr_sel == 8'hb3;
  assign mem_179_2_W0_addr = W0_addr[25:0];
  assign mem_179_2_W0_clk = W0_clk;
  assign mem_179_2_W0_data = W0_data[23:16];
  assign mem_179_2_W0_en = W0_en & W0_addr_sel == 8'hb3;
  assign mem_179_2_W0_mask = W0_mask[2];
  assign mem_179_3_R0_addr = R0_addr[25:0];
  assign mem_179_3_R0_clk = R0_clk;
  assign mem_179_3_R0_en = R0_en & R0_addr_sel == 8'hb3;
  assign mem_179_3_W0_addr = W0_addr[25:0];
  assign mem_179_3_W0_clk = W0_clk;
  assign mem_179_3_W0_data = W0_data[31:24];
  assign mem_179_3_W0_en = W0_en & W0_addr_sel == 8'hb3;
  assign mem_179_3_W0_mask = W0_mask[3];
  assign mem_179_4_R0_addr = R0_addr[25:0];
  assign mem_179_4_R0_clk = R0_clk;
  assign mem_179_4_R0_en = R0_en & R0_addr_sel == 8'hb3;
  assign mem_179_4_W0_addr = W0_addr[25:0];
  assign mem_179_4_W0_clk = W0_clk;
  assign mem_179_4_W0_data = W0_data[39:32];
  assign mem_179_4_W0_en = W0_en & W0_addr_sel == 8'hb3;
  assign mem_179_4_W0_mask = W0_mask[4];
  assign mem_179_5_R0_addr = R0_addr[25:0];
  assign mem_179_5_R0_clk = R0_clk;
  assign mem_179_5_R0_en = R0_en & R0_addr_sel == 8'hb3;
  assign mem_179_5_W0_addr = W0_addr[25:0];
  assign mem_179_5_W0_clk = W0_clk;
  assign mem_179_5_W0_data = W0_data[47:40];
  assign mem_179_5_W0_en = W0_en & W0_addr_sel == 8'hb3;
  assign mem_179_5_W0_mask = W0_mask[5];
  assign mem_179_6_R0_addr = R0_addr[25:0];
  assign mem_179_6_R0_clk = R0_clk;
  assign mem_179_6_R0_en = R0_en & R0_addr_sel == 8'hb3;
  assign mem_179_6_W0_addr = W0_addr[25:0];
  assign mem_179_6_W0_clk = W0_clk;
  assign mem_179_6_W0_data = W0_data[55:48];
  assign mem_179_6_W0_en = W0_en & W0_addr_sel == 8'hb3;
  assign mem_179_6_W0_mask = W0_mask[6];
  assign mem_179_7_R0_addr = R0_addr[25:0];
  assign mem_179_7_R0_clk = R0_clk;
  assign mem_179_7_R0_en = R0_en & R0_addr_sel == 8'hb3;
  assign mem_179_7_W0_addr = W0_addr[25:0];
  assign mem_179_7_W0_clk = W0_clk;
  assign mem_179_7_W0_data = W0_data[63:56];
  assign mem_179_7_W0_en = W0_en & W0_addr_sel == 8'hb3;
  assign mem_179_7_W0_mask = W0_mask[7];
  assign mem_180_0_R0_addr = R0_addr[25:0];
  assign mem_180_0_R0_clk = R0_clk;
  assign mem_180_0_R0_en = R0_en & R0_addr_sel == 8'hb4;
  assign mem_180_0_W0_addr = W0_addr[25:0];
  assign mem_180_0_W0_clk = W0_clk;
  assign mem_180_0_W0_data = W0_data[7:0];
  assign mem_180_0_W0_en = W0_en & W0_addr_sel == 8'hb4;
  assign mem_180_0_W0_mask = W0_mask[0];
  assign mem_180_1_R0_addr = R0_addr[25:0];
  assign mem_180_1_R0_clk = R0_clk;
  assign mem_180_1_R0_en = R0_en & R0_addr_sel == 8'hb4;
  assign mem_180_1_W0_addr = W0_addr[25:0];
  assign mem_180_1_W0_clk = W0_clk;
  assign mem_180_1_W0_data = W0_data[15:8];
  assign mem_180_1_W0_en = W0_en & W0_addr_sel == 8'hb4;
  assign mem_180_1_W0_mask = W0_mask[1];
  assign mem_180_2_R0_addr = R0_addr[25:0];
  assign mem_180_2_R0_clk = R0_clk;
  assign mem_180_2_R0_en = R0_en & R0_addr_sel == 8'hb4;
  assign mem_180_2_W0_addr = W0_addr[25:0];
  assign mem_180_2_W0_clk = W0_clk;
  assign mem_180_2_W0_data = W0_data[23:16];
  assign mem_180_2_W0_en = W0_en & W0_addr_sel == 8'hb4;
  assign mem_180_2_W0_mask = W0_mask[2];
  assign mem_180_3_R0_addr = R0_addr[25:0];
  assign mem_180_3_R0_clk = R0_clk;
  assign mem_180_3_R0_en = R0_en & R0_addr_sel == 8'hb4;
  assign mem_180_3_W0_addr = W0_addr[25:0];
  assign mem_180_3_W0_clk = W0_clk;
  assign mem_180_3_W0_data = W0_data[31:24];
  assign mem_180_3_W0_en = W0_en & W0_addr_sel == 8'hb4;
  assign mem_180_3_W0_mask = W0_mask[3];
  assign mem_180_4_R0_addr = R0_addr[25:0];
  assign mem_180_4_R0_clk = R0_clk;
  assign mem_180_4_R0_en = R0_en & R0_addr_sel == 8'hb4;
  assign mem_180_4_W0_addr = W0_addr[25:0];
  assign mem_180_4_W0_clk = W0_clk;
  assign mem_180_4_W0_data = W0_data[39:32];
  assign mem_180_4_W0_en = W0_en & W0_addr_sel == 8'hb4;
  assign mem_180_4_W0_mask = W0_mask[4];
  assign mem_180_5_R0_addr = R0_addr[25:0];
  assign mem_180_5_R0_clk = R0_clk;
  assign mem_180_5_R0_en = R0_en & R0_addr_sel == 8'hb4;
  assign mem_180_5_W0_addr = W0_addr[25:0];
  assign mem_180_5_W0_clk = W0_clk;
  assign mem_180_5_W0_data = W0_data[47:40];
  assign mem_180_5_W0_en = W0_en & W0_addr_sel == 8'hb4;
  assign mem_180_5_W0_mask = W0_mask[5];
  assign mem_180_6_R0_addr = R0_addr[25:0];
  assign mem_180_6_R0_clk = R0_clk;
  assign mem_180_6_R0_en = R0_en & R0_addr_sel == 8'hb4;
  assign mem_180_6_W0_addr = W0_addr[25:0];
  assign mem_180_6_W0_clk = W0_clk;
  assign mem_180_6_W0_data = W0_data[55:48];
  assign mem_180_6_W0_en = W0_en & W0_addr_sel == 8'hb4;
  assign mem_180_6_W0_mask = W0_mask[6];
  assign mem_180_7_R0_addr = R0_addr[25:0];
  assign mem_180_7_R0_clk = R0_clk;
  assign mem_180_7_R0_en = R0_en & R0_addr_sel == 8'hb4;
  assign mem_180_7_W0_addr = W0_addr[25:0];
  assign mem_180_7_W0_clk = W0_clk;
  assign mem_180_7_W0_data = W0_data[63:56];
  assign mem_180_7_W0_en = W0_en & W0_addr_sel == 8'hb4;
  assign mem_180_7_W0_mask = W0_mask[7];
  assign mem_181_0_R0_addr = R0_addr[25:0];
  assign mem_181_0_R0_clk = R0_clk;
  assign mem_181_0_R0_en = R0_en & R0_addr_sel == 8'hb5;
  assign mem_181_0_W0_addr = W0_addr[25:0];
  assign mem_181_0_W0_clk = W0_clk;
  assign mem_181_0_W0_data = W0_data[7:0];
  assign mem_181_0_W0_en = W0_en & W0_addr_sel == 8'hb5;
  assign mem_181_0_W0_mask = W0_mask[0];
  assign mem_181_1_R0_addr = R0_addr[25:0];
  assign mem_181_1_R0_clk = R0_clk;
  assign mem_181_1_R0_en = R0_en & R0_addr_sel == 8'hb5;
  assign mem_181_1_W0_addr = W0_addr[25:0];
  assign mem_181_1_W0_clk = W0_clk;
  assign mem_181_1_W0_data = W0_data[15:8];
  assign mem_181_1_W0_en = W0_en & W0_addr_sel == 8'hb5;
  assign mem_181_1_W0_mask = W0_mask[1];
  assign mem_181_2_R0_addr = R0_addr[25:0];
  assign mem_181_2_R0_clk = R0_clk;
  assign mem_181_2_R0_en = R0_en & R0_addr_sel == 8'hb5;
  assign mem_181_2_W0_addr = W0_addr[25:0];
  assign mem_181_2_W0_clk = W0_clk;
  assign mem_181_2_W0_data = W0_data[23:16];
  assign mem_181_2_W0_en = W0_en & W0_addr_sel == 8'hb5;
  assign mem_181_2_W0_mask = W0_mask[2];
  assign mem_181_3_R0_addr = R0_addr[25:0];
  assign mem_181_3_R0_clk = R0_clk;
  assign mem_181_3_R0_en = R0_en & R0_addr_sel == 8'hb5;
  assign mem_181_3_W0_addr = W0_addr[25:0];
  assign mem_181_3_W0_clk = W0_clk;
  assign mem_181_3_W0_data = W0_data[31:24];
  assign mem_181_3_W0_en = W0_en & W0_addr_sel == 8'hb5;
  assign mem_181_3_W0_mask = W0_mask[3];
  assign mem_181_4_R0_addr = R0_addr[25:0];
  assign mem_181_4_R0_clk = R0_clk;
  assign mem_181_4_R0_en = R0_en & R0_addr_sel == 8'hb5;
  assign mem_181_4_W0_addr = W0_addr[25:0];
  assign mem_181_4_W0_clk = W0_clk;
  assign mem_181_4_W0_data = W0_data[39:32];
  assign mem_181_4_W0_en = W0_en & W0_addr_sel == 8'hb5;
  assign mem_181_4_W0_mask = W0_mask[4];
  assign mem_181_5_R0_addr = R0_addr[25:0];
  assign mem_181_5_R0_clk = R0_clk;
  assign mem_181_5_R0_en = R0_en & R0_addr_sel == 8'hb5;
  assign mem_181_5_W0_addr = W0_addr[25:0];
  assign mem_181_5_W0_clk = W0_clk;
  assign mem_181_5_W0_data = W0_data[47:40];
  assign mem_181_5_W0_en = W0_en & W0_addr_sel == 8'hb5;
  assign mem_181_5_W0_mask = W0_mask[5];
  assign mem_181_6_R0_addr = R0_addr[25:0];
  assign mem_181_6_R0_clk = R0_clk;
  assign mem_181_6_R0_en = R0_en & R0_addr_sel == 8'hb5;
  assign mem_181_6_W0_addr = W0_addr[25:0];
  assign mem_181_6_W0_clk = W0_clk;
  assign mem_181_6_W0_data = W0_data[55:48];
  assign mem_181_6_W0_en = W0_en & W0_addr_sel == 8'hb5;
  assign mem_181_6_W0_mask = W0_mask[6];
  assign mem_181_7_R0_addr = R0_addr[25:0];
  assign mem_181_7_R0_clk = R0_clk;
  assign mem_181_7_R0_en = R0_en & R0_addr_sel == 8'hb5;
  assign mem_181_7_W0_addr = W0_addr[25:0];
  assign mem_181_7_W0_clk = W0_clk;
  assign mem_181_7_W0_data = W0_data[63:56];
  assign mem_181_7_W0_en = W0_en & W0_addr_sel == 8'hb5;
  assign mem_181_7_W0_mask = W0_mask[7];
  assign mem_182_0_R0_addr = R0_addr[25:0];
  assign mem_182_0_R0_clk = R0_clk;
  assign mem_182_0_R0_en = R0_en & R0_addr_sel == 8'hb6;
  assign mem_182_0_W0_addr = W0_addr[25:0];
  assign mem_182_0_W0_clk = W0_clk;
  assign mem_182_0_W0_data = W0_data[7:0];
  assign mem_182_0_W0_en = W0_en & W0_addr_sel == 8'hb6;
  assign mem_182_0_W0_mask = W0_mask[0];
  assign mem_182_1_R0_addr = R0_addr[25:0];
  assign mem_182_1_R0_clk = R0_clk;
  assign mem_182_1_R0_en = R0_en & R0_addr_sel == 8'hb6;
  assign mem_182_1_W0_addr = W0_addr[25:0];
  assign mem_182_1_W0_clk = W0_clk;
  assign mem_182_1_W0_data = W0_data[15:8];
  assign mem_182_1_W0_en = W0_en & W0_addr_sel == 8'hb6;
  assign mem_182_1_W0_mask = W0_mask[1];
  assign mem_182_2_R0_addr = R0_addr[25:0];
  assign mem_182_2_R0_clk = R0_clk;
  assign mem_182_2_R0_en = R0_en & R0_addr_sel == 8'hb6;
  assign mem_182_2_W0_addr = W0_addr[25:0];
  assign mem_182_2_W0_clk = W0_clk;
  assign mem_182_2_W0_data = W0_data[23:16];
  assign mem_182_2_W0_en = W0_en & W0_addr_sel == 8'hb6;
  assign mem_182_2_W0_mask = W0_mask[2];
  assign mem_182_3_R0_addr = R0_addr[25:0];
  assign mem_182_3_R0_clk = R0_clk;
  assign mem_182_3_R0_en = R0_en & R0_addr_sel == 8'hb6;
  assign mem_182_3_W0_addr = W0_addr[25:0];
  assign mem_182_3_W0_clk = W0_clk;
  assign mem_182_3_W0_data = W0_data[31:24];
  assign mem_182_3_W0_en = W0_en & W0_addr_sel == 8'hb6;
  assign mem_182_3_W0_mask = W0_mask[3];
  assign mem_182_4_R0_addr = R0_addr[25:0];
  assign mem_182_4_R0_clk = R0_clk;
  assign mem_182_4_R0_en = R0_en & R0_addr_sel == 8'hb6;
  assign mem_182_4_W0_addr = W0_addr[25:0];
  assign mem_182_4_W0_clk = W0_clk;
  assign mem_182_4_W0_data = W0_data[39:32];
  assign mem_182_4_W0_en = W0_en & W0_addr_sel == 8'hb6;
  assign mem_182_4_W0_mask = W0_mask[4];
  assign mem_182_5_R0_addr = R0_addr[25:0];
  assign mem_182_5_R0_clk = R0_clk;
  assign mem_182_5_R0_en = R0_en & R0_addr_sel == 8'hb6;
  assign mem_182_5_W0_addr = W0_addr[25:0];
  assign mem_182_5_W0_clk = W0_clk;
  assign mem_182_5_W0_data = W0_data[47:40];
  assign mem_182_5_W0_en = W0_en & W0_addr_sel == 8'hb6;
  assign mem_182_5_W0_mask = W0_mask[5];
  assign mem_182_6_R0_addr = R0_addr[25:0];
  assign mem_182_6_R0_clk = R0_clk;
  assign mem_182_6_R0_en = R0_en & R0_addr_sel == 8'hb6;
  assign mem_182_6_W0_addr = W0_addr[25:0];
  assign mem_182_6_W0_clk = W0_clk;
  assign mem_182_6_W0_data = W0_data[55:48];
  assign mem_182_6_W0_en = W0_en & W0_addr_sel == 8'hb6;
  assign mem_182_6_W0_mask = W0_mask[6];
  assign mem_182_7_R0_addr = R0_addr[25:0];
  assign mem_182_7_R0_clk = R0_clk;
  assign mem_182_7_R0_en = R0_en & R0_addr_sel == 8'hb6;
  assign mem_182_7_W0_addr = W0_addr[25:0];
  assign mem_182_7_W0_clk = W0_clk;
  assign mem_182_7_W0_data = W0_data[63:56];
  assign mem_182_7_W0_en = W0_en & W0_addr_sel == 8'hb6;
  assign mem_182_7_W0_mask = W0_mask[7];
  assign mem_183_0_R0_addr = R0_addr[25:0];
  assign mem_183_0_R0_clk = R0_clk;
  assign mem_183_0_R0_en = R0_en & R0_addr_sel == 8'hb7;
  assign mem_183_0_W0_addr = W0_addr[25:0];
  assign mem_183_0_W0_clk = W0_clk;
  assign mem_183_0_W0_data = W0_data[7:0];
  assign mem_183_0_W0_en = W0_en & W0_addr_sel == 8'hb7;
  assign mem_183_0_W0_mask = W0_mask[0];
  assign mem_183_1_R0_addr = R0_addr[25:0];
  assign mem_183_1_R0_clk = R0_clk;
  assign mem_183_1_R0_en = R0_en & R0_addr_sel == 8'hb7;
  assign mem_183_1_W0_addr = W0_addr[25:0];
  assign mem_183_1_W0_clk = W0_clk;
  assign mem_183_1_W0_data = W0_data[15:8];
  assign mem_183_1_W0_en = W0_en & W0_addr_sel == 8'hb7;
  assign mem_183_1_W0_mask = W0_mask[1];
  assign mem_183_2_R0_addr = R0_addr[25:0];
  assign mem_183_2_R0_clk = R0_clk;
  assign mem_183_2_R0_en = R0_en & R0_addr_sel == 8'hb7;
  assign mem_183_2_W0_addr = W0_addr[25:0];
  assign mem_183_2_W0_clk = W0_clk;
  assign mem_183_2_W0_data = W0_data[23:16];
  assign mem_183_2_W0_en = W0_en & W0_addr_sel == 8'hb7;
  assign mem_183_2_W0_mask = W0_mask[2];
  assign mem_183_3_R0_addr = R0_addr[25:0];
  assign mem_183_3_R0_clk = R0_clk;
  assign mem_183_3_R0_en = R0_en & R0_addr_sel == 8'hb7;
  assign mem_183_3_W0_addr = W0_addr[25:0];
  assign mem_183_3_W0_clk = W0_clk;
  assign mem_183_3_W0_data = W0_data[31:24];
  assign mem_183_3_W0_en = W0_en & W0_addr_sel == 8'hb7;
  assign mem_183_3_W0_mask = W0_mask[3];
  assign mem_183_4_R0_addr = R0_addr[25:0];
  assign mem_183_4_R0_clk = R0_clk;
  assign mem_183_4_R0_en = R0_en & R0_addr_sel == 8'hb7;
  assign mem_183_4_W0_addr = W0_addr[25:0];
  assign mem_183_4_W0_clk = W0_clk;
  assign mem_183_4_W0_data = W0_data[39:32];
  assign mem_183_4_W0_en = W0_en & W0_addr_sel == 8'hb7;
  assign mem_183_4_W0_mask = W0_mask[4];
  assign mem_183_5_R0_addr = R0_addr[25:0];
  assign mem_183_5_R0_clk = R0_clk;
  assign mem_183_5_R0_en = R0_en & R0_addr_sel == 8'hb7;
  assign mem_183_5_W0_addr = W0_addr[25:0];
  assign mem_183_5_W0_clk = W0_clk;
  assign mem_183_5_W0_data = W0_data[47:40];
  assign mem_183_5_W0_en = W0_en & W0_addr_sel == 8'hb7;
  assign mem_183_5_W0_mask = W0_mask[5];
  assign mem_183_6_R0_addr = R0_addr[25:0];
  assign mem_183_6_R0_clk = R0_clk;
  assign mem_183_6_R0_en = R0_en & R0_addr_sel == 8'hb7;
  assign mem_183_6_W0_addr = W0_addr[25:0];
  assign mem_183_6_W0_clk = W0_clk;
  assign mem_183_6_W0_data = W0_data[55:48];
  assign mem_183_6_W0_en = W0_en & W0_addr_sel == 8'hb7;
  assign mem_183_6_W0_mask = W0_mask[6];
  assign mem_183_7_R0_addr = R0_addr[25:0];
  assign mem_183_7_R0_clk = R0_clk;
  assign mem_183_7_R0_en = R0_en & R0_addr_sel == 8'hb7;
  assign mem_183_7_W0_addr = W0_addr[25:0];
  assign mem_183_7_W0_clk = W0_clk;
  assign mem_183_7_W0_data = W0_data[63:56];
  assign mem_183_7_W0_en = W0_en & W0_addr_sel == 8'hb7;
  assign mem_183_7_W0_mask = W0_mask[7];
  assign mem_184_0_R0_addr = R0_addr[25:0];
  assign mem_184_0_R0_clk = R0_clk;
  assign mem_184_0_R0_en = R0_en & R0_addr_sel == 8'hb8;
  assign mem_184_0_W0_addr = W0_addr[25:0];
  assign mem_184_0_W0_clk = W0_clk;
  assign mem_184_0_W0_data = W0_data[7:0];
  assign mem_184_0_W0_en = W0_en & W0_addr_sel == 8'hb8;
  assign mem_184_0_W0_mask = W0_mask[0];
  assign mem_184_1_R0_addr = R0_addr[25:0];
  assign mem_184_1_R0_clk = R0_clk;
  assign mem_184_1_R0_en = R0_en & R0_addr_sel == 8'hb8;
  assign mem_184_1_W0_addr = W0_addr[25:0];
  assign mem_184_1_W0_clk = W0_clk;
  assign mem_184_1_W0_data = W0_data[15:8];
  assign mem_184_1_W0_en = W0_en & W0_addr_sel == 8'hb8;
  assign mem_184_1_W0_mask = W0_mask[1];
  assign mem_184_2_R0_addr = R0_addr[25:0];
  assign mem_184_2_R0_clk = R0_clk;
  assign mem_184_2_R0_en = R0_en & R0_addr_sel == 8'hb8;
  assign mem_184_2_W0_addr = W0_addr[25:0];
  assign mem_184_2_W0_clk = W0_clk;
  assign mem_184_2_W0_data = W0_data[23:16];
  assign mem_184_2_W0_en = W0_en & W0_addr_sel == 8'hb8;
  assign mem_184_2_W0_mask = W0_mask[2];
  assign mem_184_3_R0_addr = R0_addr[25:0];
  assign mem_184_3_R0_clk = R0_clk;
  assign mem_184_3_R0_en = R0_en & R0_addr_sel == 8'hb8;
  assign mem_184_3_W0_addr = W0_addr[25:0];
  assign mem_184_3_W0_clk = W0_clk;
  assign mem_184_3_W0_data = W0_data[31:24];
  assign mem_184_3_W0_en = W0_en & W0_addr_sel == 8'hb8;
  assign mem_184_3_W0_mask = W0_mask[3];
  assign mem_184_4_R0_addr = R0_addr[25:0];
  assign mem_184_4_R0_clk = R0_clk;
  assign mem_184_4_R0_en = R0_en & R0_addr_sel == 8'hb8;
  assign mem_184_4_W0_addr = W0_addr[25:0];
  assign mem_184_4_W0_clk = W0_clk;
  assign mem_184_4_W0_data = W0_data[39:32];
  assign mem_184_4_W0_en = W0_en & W0_addr_sel == 8'hb8;
  assign mem_184_4_W0_mask = W0_mask[4];
  assign mem_184_5_R0_addr = R0_addr[25:0];
  assign mem_184_5_R0_clk = R0_clk;
  assign mem_184_5_R0_en = R0_en & R0_addr_sel == 8'hb8;
  assign mem_184_5_W0_addr = W0_addr[25:0];
  assign mem_184_5_W0_clk = W0_clk;
  assign mem_184_5_W0_data = W0_data[47:40];
  assign mem_184_5_W0_en = W0_en & W0_addr_sel == 8'hb8;
  assign mem_184_5_W0_mask = W0_mask[5];
  assign mem_184_6_R0_addr = R0_addr[25:0];
  assign mem_184_6_R0_clk = R0_clk;
  assign mem_184_6_R0_en = R0_en & R0_addr_sel == 8'hb8;
  assign mem_184_6_W0_addr = W0_addr[25:0];
  assign mem_184_6_W0_clk = W0_clk;
  assign mem_184_6_W0_data = W0_data[55:48];
  assign mem_184_6_W0_en = W0_en & W0_addr_sel == 8'hb8;
  assign mem_184_6_W0_mask = W0_mask[6];
  assign mem_184_7_R0_addr = R0_addr[25:0];
  assign mem_184_7_R0_clk = R0_clk;
  assign mem_184_7_R0_en = R0_en & R0_addr_sel == 8'hb8;
  assign mem_184_7_W0_addr = W0_addr[25:0];
  assign mem_184_7_W0_clk = W0_clk;
  assign mem_184_7_W0_data = W0_data[63:56];
  assign mem_184_7_W0_en = W0_en & W0_addr_sel == 8'hb8;
  assign mem_184_7_W0_mask = W0_mask[7];
  assign mem_185_0_R0_addr = R0_addr[25:0];
  assign mem_185_0_R0_clk = R0_clk;
  assign mem_185_0_R0_en = R0_en & R0_addr_sel == 8'hb9;
  assign mem_185_0_W0_addr = W0_addr[25:0];
  assign mem_185_0_W0_clk = W0_clk;
  assign mem_185_0_W0_data = W0_data[7:0];
  assign mem_185_0_W0_en = W0_en & W0_addr_sel == 8'hb9;
  assign mem_185_0_W0_mask = W0_mask[0];
  assign mem_185_1_R0_addr = R0_addr[25:0];
  assign mem_185_1_R0_clk = R0_clk;
  assign mem_185_1_R0_en = R0_en & R0_addr_sel == 8'hb9;
  assign mem_185_1_W0_addr = W0_addr[25:0];
  assign mem_185_1_W0_clk = W0_clk;
  assign mem_185_1_W0_data = W0_data[15:8];
  assign mem_185_1_W0_en = W0_en & W0_addr_sel == 8'hb9;
  assign mem_185_1_W0_mask = W0_mask[1];
  assign mem_185_2_R0_addr = R0_addr[25:0];
  assign mem_185_2_R0_clk = R0_clk;
  assign mem_185_2_R0_en = R0_en & R0_addr_sel == 8'hb9;
  assign mem_185_2_W0_addr = W0_addr[25:0];
  assign mem_185_2_W0_clk = W0_clk;
  assign mem_185_2_W0_data = W0_data[23:16];
  assign mem_185_2_W0_en = W0_en & W0_addr_sel == 8'hb9;
  assign mem_185_2_W0_mask = W0_mask[2];
  assign mem_185_3_R0_addr = R0_addr[25:0];
  assign mem_185_3_R0_clk = R0_clk;
  assign mem_185_3_R0_en = R0_en & R0_addr_sel == 8'hb9;
  assign mem_185_3_W0_addr = W0_addr[25:0];
  assign mem_185_3_W0_clk = W0_clk;
  assign mem_185_3_W0_data = W0_data[31:24];
  assign mem_185_3_W0_en = W0_en & W0_addr_sel == 8'hb9;
  assign mem_185_3_W0_mask = W0_mask[3];
  assign mem_185_4_R0_addr = R0_addr[25:0];
  assign mem_185_4_R0_clk = R0_clk;
  assign mem_185_4_R0_en = R0_en & R0_addr_sel == 8'hb9;
  assign mem_185_4_W0_addr = W0_addr[25:0];
  assign mem_185_4_W0_clk = W0_clk;
  assign mem_185_4_W0_data = W0_data[39:32];
  assign mem_185_4_W0_en = W0_en & W0_addr_sel == 8'hb9;
  assign mem_185_4_W0_mask = W0_mask[4];
  assign mem_185_5_R0_addr = R0_addr[25:0];
  assign mem_185_5_R0_clk = R0_clk;
  assign mem_185_5_R0_en = R0_en & R0_addr_sel == 8'hb9;
  assign mem_185_5_W0_addr = W0_addr[25:0];
  assign mem_185_5_W0_clk = W0_clk;
  assign mem_185_5_W0_data = W0_data[47:40];
  assign mem_185_5_W0_en = W0_en & W0_addr_sel == 8'hb9;
  assign mem_185_5_W0_mask = W0_mask[5];
  assign mem_185_6_R0_addr = R0_addr[25:0];
  assign mem_185_6_R0_clk = R0_clk;
  assign mem_185_6_R0_en = R0_en & R0_addr_sel == 8'hb9;
  assign mem_185_6_W0_addr = W0_addr[25:0];
  assign mem_185_6_W0_clk = W0_clk;
  assign mem_185_6_W0_data = W0_data[55:48];
  assign mem_185_6_W0_en = W0_en & W0_addr_sel == 8'hb9;
  assign mem_185_6_W0_mask = W0_mask[6];
  assign mem_185_7_R0_addr = R0_addr[25:0];
  assign mem_185_7_R0_clk = R0_clk;
  assign mem_185_7_R0_en = R0_en & R0_addr_sel == 8'hb9;
  assign mem_185_7_W0_addr = W0_addr[25:0];
  assign mem_185_7_W0_clk = W0_clk;
  assign mem_185_7_W0_data = W0_data[63:56];
  assign mem_185_7_W0_en = W0_en & W0_addr_sel == 8'hb9;
  assign mem_185_7_W0_mask = W0_mask[7];
  assign mem_186_0_R0_addr = R0_addr[25:0];
  assign mem_186_0_R0_clk = R0_clk;
  assign mem_186_0_R0_en = R0_en & R0_addr_sel == 8'hba;
  assign mem_186_0_W0_addr = W0_addr[25:0];
  assign mem_186_0_W0_clk = W0_clk;
  assign mem_186_0_W0_data = W0_data[7:0];
  assign mem_186_0_W0_en = W0_en & W0_addr_sel == 8'hba;
  assign mem_186_0_W0_mask = W0_mask[0];
  assign mem_186_1_R0_addr = R0_addr[25:0];
  assign mem_186_1_R0_clk = R0_clk;
  assign mem_186_1_R0_en = R0_en & R0_addr_sel == 8'hba;
  assign mem_186_1_W0_addr = W0_addr[25:0];
  assign mem_186_1_W0_clk = W0_clk;
  assign mem_186_1_W0_data = W0_data[15:8];
  assign mem_186_1_W0_en = W0_en & W0_addr_sel == 8'hba;
  assign mem_186_1_W0_mask = W0_mask[1];
  assign mem_186_2_R0_addr = R0_addr[25:0];
  assign mem_186_2_R0_clk = R0_clk;
  assign mem_186_2_R0_en = R0_en & R0_addr_sel == 8'hba;
  assign mem_186_2_W0_addr = W0_addr[25:0];
  assign mem_186_2_W0_clk = W0_clk;
  assign mem_186_2_W0_data = W0_data[23:16];
  assign mem_186_2_W0_en = W0_en & W0_addr_sel == 8'hba;
  assign mem_186_2_W0_mask = W0_mask[2];
  assign mem_186_3_R0_addr = R0_addr[25:0];
  assign mem_186_3_R0_clk = R0_clk;
  assign mem_186_3_R0_en = R0_en & R0_addr_sel == 8'hba;
  assign mem_186_3_W0_addr = W0_addr[25:0];
  assign mem_186_3_W0_clk = W0_clk;
  assign mem_186_3_W0_data = W0_data[31:24];
  assign mem_186_3_W0_en = W0_en & W0_addr_sel == 8'hba;
  assign mem_186_3_W0_mask = W0_mask[3];
  assign mem_186_4_R0_addr = R0_addr[25:0];
  assign mem_186_4_R0_clk = R0_clk;
  assign mem_186_4_R0_en = R0_en & R0_addr_sel == 8'hba;
  assign mem_186_4_W0_addr = W0_addr[25:0];
  assign mem_186_4_W0_clk = W0_clk;
  assign mem_186_4_W0_data = W0_data[39:32];
  assign mem_186_4_W0_en = W0_en & W0_addr_sel == 8'hba;
  assign mem_186_4_W0_mask = W0_mask[4];
  assign mem_186_5_R0_addr = R0_addr[25:0];
  assign mem_186_5_R0_clk = R0_clk;
  assign mem_186_5_R0_en = R0_en & R0_addr_sel == 8'hba;
  assign mem_186_5_W0_addr = W0_addr[25:0];
  assign mem_186_5_W0_clk = W0_clk;
  assign mem_186_5_W0_data = W0_data[47:40];
  assign mem_186_5_W0_en = W0_en & W0_addr_sel == 8'hba;
  assign mem_186_5_W0_mask = W0_mask[5];
  assign mem_186_6_R0_addr = R0_addr[25:0];
  assign mem_186_6_R0_clk = R0_clk;
  assign mem_186_6_R0_en = R0_en & R0_addr_sel == 8'hba;
  assign mem_186_6_W0_addr = W0_addr[25:0];
  assign mem_186_6_W0_clk = W0_clk;
  assign mem_186_6_W0_data = W0_data[55:48];
  assign mem_186_6_W0_en = W0_en & W0_addr_sel == 8'hba;
  assign mem_186_6_W0_mask = W0_mask[6];
  assign mem_186_7_R0_addr = R0_addr[25:0];
  assign mem_186_7_R0_clk = R0_clk;
  assign mem_186_7_R0_en = R0_en & R0_addr_sel == 8'hba;
  assign mem_186_7_W0_addr = W0_addr[25:0];
  assign mem_186_7_W0_clk = W0_clk;
  assign mem_186_7_W0_data = W0_data[63:56];
  assign mem_186_7_W0_en = W0_en & W0_addr_sel == 8'hba;
  assign mem_186_7_W0_mask = W0_mask[7];
  assign mem_187_0_R0_addr = R0_addr[25:0];
  assign mem_187_0_R0_clk = R0_clk;
  assign mem_187_0_R0_en = R0_en & R0_addr_sel == 8'hbb;
  assign mem_187_0_W0_addr = W0_addr[25:0];
  assign mem_187_0_W0_clk = W0_clk;
  assign mem_187_0_W0_data = W0_data[7:0];
  assign mem_187_0_W0_en = W0_en & W0_addr_sel == 8'hbb;
  assign mem_187_0_W0_mask = W0_mask[0];
  assign mem_187_1_R0_addr = R0_addr[25:0];
  assign mem_187_1_R0_clk = R0_clk;
  assign mem_187_1_R0_en = R0_en & R0_addr_sel == 8'hbb;
  assign mem_187_1_W0_addr = W0_addr[25:0];
  assign mem_187_1_W0_clk = W0_clk;
  assign mem_187_1_W0_data = W0_data[15:8];
  assign mem_187_1_W0_en = W0_en & W0_addr_sel == 8'hbb;
  assign mem_187_1_W0_mask = W0_mask[1];
  assign mem_187_2_R0_addr = R0_addr[25:0];
  assign mem_187_2_R0_clk = R0_clk;
  assign mem_187_2_R0_en = R0_en & R0_addr_sel == 8'hbb;
  assign mem_187_2_W0_addr = W0_addr[25:0];
  assign mem_187_2_W0_clk = W0_clk;
  assign mem_187_2_W0_data = W0_data[23:16];
  assign mem_187_2_W0_en = W0_en & W0_addr_sel == 8'hbb;
  assign mem_187_2_W0_mask = W0_mask[2];
  assign mem_187_3_R0_addr = R0_addr[25:0];
  assign mem_187_3_R0_clk = R0_clk;
  assign mem_187_3_R0_en = R0_en & R0_addr_sel == 8'hbb;
  assign mem_187_3_W0_addr = W0_addr[25:0];
  assign mem_187_3_W0_clk = W0_clk;
  assign mem_187_3_W0_data = W0_data[31:24];
  assign mem_187_3_W0_en = W0_en & W0_addr_sel == 8'hbb;
  assign mem_187_3_W0_mask = W0_mask[3];
  assign mem_187_4_R0_addr = R0_addr[25:0];
  assign mem_187_4_R0_clk = R0_clk;
  assign mem_187_4_R0_en = R0_en & R0_addr_sel == 8'hbb;
  assign mem_187_4_W0_addr = W0_addr[25:0];
  assign mem_187_4_W0_clk = W0_clk;
  assign mem_187_4_W0_data = W0_data[39:32];
  assign mem_187_4_W0_en = W0_en & W0_addr_sel == 8'hbb;
  assign mem_187_4_W0_mask = W0_mask[4];
  assign mem_187_5_R0_addr = R0_addr[25:0];
  assign mem_187_5_R0_clk = R0_clk;
  assign mem_187_5_R0_en = R0_en & R0_addr_sel == 8'hbb;
  assign mem_187_5_W0_addr = W0_addr[25:0];
  assign mem_187_5_W0_clk = W0_clk;
  assign mem_187_5_W0_data = W0_data[47:40];
  assign mem_187_5_W0_en = W0_en & W0_addr_sel == 8'hbb;
  assign mem_187_5_W0_mask = W0_mask[5];
  assign mem_187_6_R0_addr = R0_addr[25:0];
  assign mem_187_6_R0_clk = R0_clk;
  assign mem_187_6_R0_en = R0_en & R0_addr_sel == 8'hbb;
  assign mem_187_6_W0_addr = W0_addr[25:0];
  assign mem_187_6_W0_clk = W0_clk;
  assign mem_187_6_W0_data = W0_data[55:48];
  assign mem_187_6_W0_en = W0_en & W0_addr_sel == 8'hbb;
  assign mem_187_6_W0_mask = W0_mask[6];
  assign mem_187_7_R0_addr = R0_addr[25:0];
  assign mem_187_7_R0_clk = R0_clk;
  assign mem_187_7_R0_en = R0_en & R0_addr_sel == 8'hbb;
  assign mem_187_7_W0_addr = W0_addr[25:0];
  assign mem_187_7_W0_clk = W0_clk;
  assign mem_187_7_W0_data = W0_data[63:56];
  assign mem_187_7_W0_en = W0_en & W0_addr_sel == 8'hbb;
  assign mem_187_7_W0_mask = W0_mask[7];
  assign mem_188_0_R0_addr = R0_addr[25:0];
  assign mem_188_0_R0_clk = R0_clk;
  assign mem_188_0_R0_en = R0_en & R0_addr_sel == 8'hbc;
  assign mem_188_0_W0_addr = W0_addr[25:0];
  assign mem_188_0_W0_clk = W0_clk;
  assign mem_188_0_W0_data = W0_data[7:0];
  assign mem_188_0_W0_en = W0_en & W0_addr_sel == 8'hbc;
  assign mem_188_0_W0_mask = W0_mask[0];
  assign mem_188_1_R0_addr = R0_addr[25:0];
  assign mem_188_1_R0_clk = R0_clk;
  assign mem_188_1_R0_en = R0_en & R0_addr_sel == 8'hbc;
  assign mem_188_1_W0_addr = W0_addr[25:0];
  assign mem_188_1_W0_clk = W0_clk;
  assign mem_188_1_W0_data = W0_data[15:8];
  assign mem_188_1_W0_en = W0_en & W0_addr_sel == 8'hbc;
  assign mem_188_1_W0_mask = W0_mask[1];
  assign mem_188_2_R0_addr = R0_addr[25:0];
  assign mem_188_2_R0_clk = R0_clk;
  assign mem_188_2_R0_en = R0_en & R0_addr_sel == 8'hbc;
  assign mem_188_2_W0_addr = W0_addr[25:0];
  assign mem_188_2_W0_clk = W0_clk;
  assign mem_188_2_W0_data = W0_data[23:16];
  assign mem_188_2_W0_en = W0_en & W0_addr_sel == 8'hbc;
  assign mem_188_2_W0_mask = W0_mask[2];
  assign mem_188_3_R0_addr = R0_addr[25:0];
  assign mem_188_3_R0_clk = R0_clk;
  assign mem_188_3_R0_en = R0_en & R0_addr_sel == 8'hbc;
  assign mem_188_3_W0_addr = W0_addr[25:0];
  assign mem_188_3_W0_clk = W0_clk;
  assign mem_188_3_W0_data = W0_data[31:24];
  assign mem_188_3_W0_en = W0_en & W0_addr_sel == 8'hbc;
  assign mem_188_3_W0_mask = W0_mask[3];
  assign mem_188_4_R0_addr = R0_addr[25:0];
  assign mem_188_4_R0_clk = R0_clk;
  assign mem_188_4_R0_en = R0_en & R0_addr_sel == 8'hbc;
  assign mem_188_4_W0_addr = W0_addr[25:0];
  assign mem_188_4_W0_clk = W0_clk;
  assign mem_188_4_W0_data = W0_data[39:32];
  assign mem_188_4_W0_en = W0_en & W0_addr_sel == 8'hbc;
  assign mem_188_4_W0_mask = W0_mask[4];
  assign mem_188_5_R0_addr = R0_addr[25:0];
  assign mem_188_5_R0_clk = R0_clk;
  assign mem_188_5_R0_en = R0_en & R0_addr_sel == 8'hbc;
  assign mem_188_5_W0_addr = W0_addr[25:0];
  assign mem_188_5_W0_clk = W0_clk;
  assign mem_188_5_W0_data = W0_data[47:40];
  assign mem_188_5_W0_en = W0_en & W0_addr_sel == 8'hbc;
  assign mem_188_5_W0_mask = W0_mask[5];
  assign mem_188_6_R0_addr = R0_addr[25:0];
  assign mem_188_6_R0_clk = R0_clk;
  assign mem_188_6_R0_en = R0_en & R0_addr_sel == 8'hbc;
  assign mem_188_6_W0_addr = W0_addr[25:0];
  assign mem_188_6_W0_clk = W0_clk;
  assign mem_188_6_W0_data = W0_data[55:48];
  assign mem_188_6_W0_en = W0_en & W0_addr_sel == 8'hbc;
  assign mem_188_6_W0_mask = W0_mask[6];
  assign mem_188_7_R0_addr = R0_addr[25:0];
  assign mem_188_7_R0_clk = R0_clk;
  assign mem_188_7_R0_en = R0_en & R0_addr_sel == 8'hbc;
  assign mem_188_7_W0_addr = W0_addr[25:0];
  assign mem_188_7_W0_clk = W0_clk;
  assign mem_188_7_W0_data = W0_data[63:56];
  assign mem_188_7_W0_en = W0_en & W0_addr_sel == 8'hbc;
  assign mem_188_7_W0_mask = W0_mask[7];
  assign mem_189_0_R0_addr = R0_addr[25:0];
  assign mem_189_0_R0_clk = R0_clk;
  assign mem_189_0_R0_en = R0_en & R0_addr_sel == 8'hbd;
  assign mem_189_0_W0_addr = W0_addr[25:0];
  assign mem_189_0_W0_clk = W0_clk;
  assign mem_189_0_W0_data = W0_data[7:0];
  assign mem_189_0_W0_en = W0_en & W0_addr_sel == 8'hbd;
  assign mem_189_0_W0_mask = W0_mask[0];
  assign mem_189_1_R0_addr = R0_addr[25:0];
  assign mem_189_1_R0_clk = R0_clk;
  assign mem_189_1_R0_en = R0_en & R0_addr_sel == 8'hbd;
  assign mem_189_1_W0_addr = W0_addr[25:0];
  assign mem_189_1_W0_clk = W0_clk;
  assign mem_189_1_W0_data = W0_data[15:8];
  assign mem_189_1_W0_en = W0_en & W0_addr_sel == 8'hbd;
  assign mem_189_1_W0_mask = W0_mask[1];
  assign mem_189_2_R0_addr = R0_addr[25:0];
  assign mem_189_2_R0_clk = R0_clk;
  assign mem_189_2_R0_en = R0_en & R0_addr_sel == 8'hbd;
  assign mem_189_2_W0_addr = W0_addr[25:0];
  assign mem_189_2_W0_clk = W0_clk;
  assign mem_189_2_W0_data = W0_data[23:16];
  assign mem_189_2_W0_en = W0_en & W0_addr_sel == 8'hbd;
  assign mem_189_2_W0_mask = W0_mask[2];
  assign mem_189_3_R0_addr = R0_addr[25:0];
  assign mem_189_3_R0_clk = R0_clk;
  assign mem_189_3_R0_en = R0_en & R0_addr_sel == 8'hbd;
  assign mem_189_3_W0_addr = W0_addr[25:0];
  assign mem_189_3_W0_clk = W0_clk;
  assign mem_189_3_W0_data = W0_data[31:24];
  assign mem_189_3_W0_en = W0_en & W0_addr_sel == 8'hbd;
  assign mem_189_3_W0_mask = W0_mask[3];
  assign mem_189_4_R0_addr = R0_addr[25:0];
  assign mem_189_4_R0_clk = R0_clk;
  assign mem_189_4_R0_en = R0_en & R0_addr_sel == 8'hbd;
  assign mem_189_4_W0_addr = W0_addr[25:0];
  assign mem_189_4_W0_clk = W0_clk;
  assign mem_189_4_W0_data = W0_data[39:32];
  assign mem_189_4_W0_en = W0_en & W0_addr_sel == 8'hbd;
  assign mem_189_4_W0_mask = W0_mask[4];
  assign mem_189_5_R0_addr = R0_addr[25:0];
  assign mem_189_5_R0_clk = R0_clk;
  assign mem_189_5_R0_en = R0_en & R0_addr_sel == 8'hbd;
  assign mem_189_5_W0_addr = W0_addr[25:0];
  assign mem_189_5_W0_clk = W0_clk;
  assign mem_189_5_W0_data = W0_data[47:40];
  assign mem_189_5_W0_en = W0_en & W0_addr_sel == 8'hbd;
  assign mem_189_5_W0_mask = W0_mask[5];
  assign mem_189_6_R0_addr = R0_addr[25:0];
  assign mem_189_6_R0_clk = R0_clk;
  assign mem_189_6_R0_en = R0_en & R0_addr_sel == 8'hbd;
  assign mem_189_6_W0_addr = W0_addr[25:0];
  assign mem_189_6_W0_clk = W0_clk;
  assign mem_189_6_W0_data = W0_data[55:48];
  assign mem_189_6_W0_en = W0_en & W0_addr_sel == 8'hbd;
  assign mem_189_6_W0_mask = W0_mask[6];
  assign mem_189_7_R0_addr = R0_addr[25:0];
  assign mem_189_7_R0_clk = R0_clk;
  assign mem_189_7_R0_en = R0_en & R0_addr_sel == 8'hbd;
  assign mem_189_7_W0_addr = W0_addr[25:0];
  assign mem_189_7_W0_clk = W0_clk;
  assign mem_189_7_W0_data = W0_data[63:56];
  assign mem_189_7_W0_en = W0_en & W0_addr_sel == 8'hbd;
  assign mem_189_7_W0_mask = W0_mask[7];
  assign mem_190_0_R0_addr = R0_addr[25:0];
  assign mem_190_0_R0_clk = R0_clk;
  assign mem_190_0_R0_en = R0_en & R0_addr_sel == 8'hbe;
  assign mem_190_0_W0_addr = W0_addr[25:0];
  assign mem_190_0_W0_clk = W0_clk;
  assign mem_190_0_W0_data = W0_data[7:0];
  assign mem_190_0_W0_en = W0_en & W0_addr_sel == 8'hbe;
  assign mem_190_0_W0_mask = W0_mask[0];
  assign mem_190_1_R0_addr = R0_addr[25:0];
  assign mem_190_1_R0_clk = R0_clk;
  assign mem_190_1_R0_en = R0_en & R0_addr_sel == 8'hbe;
  assign mem_190_1_W0_addr = W0_addr[25:0];
  assign mem_190_1_W0_clk = W0_clk;
  assign mem_190_1_W0_data = W0_data[15:8];
  assign mem_190_1_W0_en = W0_en & W0_addr_sel == 8'hbe;
  assign mem_190_1_W0_mask = W0_mask[1];
  assign mem_190_2_R0_addr = R0_addr[25:0];
  assign mem_190_2_R0_clk = R0_clk;
  assign mem_190_2_R0_en = R0_en & R0_addr_sel == 8'hbe;
  assign mem_190_2_W0_addr = W0_addr[25:0];
  assign mem_190_2_W0_clk = W0_clk;
  assign mem_190_2_W0_data = W0_data[23:16];
  assign mem_190_2_W0_en = W0_en & W0_addr_sel == 8'hbe;
  assign mem_190_2_W0_mask = W0_mask[2];
  assign mem_190_3_R0_addr = R0_addr[25:0];
  assign mem_190_3_R0_clk = R0_clk;
  assign mem_190_3_R0_en = R0_en & R0_addr_sel == 8'hbe;
  assign mem_190_3_W0_addr = W0_addr[25:0];
  assign mem_190_3_W0_clk = W0_clk;
  assign mem_190_3_W0_data = W0_data[31:24];
  assign mem_190_3_W0_en = W0_en & W0_addr_sel == 8'hbe;
  assign mem_190_3_W0_mask = W0_mask[3];
  assign mem_190_4_R0_addr = R0_addr[25:0];
  assign mem_190_4_R0_clk = R0_clk;
  assign mem_190_4_R0_en = R0_en & R0_addr_sel == 8'hbe;
  assign mem_190_4_W0_addr = W0_addr[25:0];
  assign mem_190_4_W0_clk = W0_clk;
  assign mem_190_4_W0_data = W0_data[39:32];
  assign mem_190_4_W0_en = W0_en & W0_addr_sel == 8'hbe;
  assign mem_190_4_W0_mask = W0_mask[4];
  assign mem_190_5_R0_addr = R0_addr[25:0];
  assign mem_190_5_R0_clk = R0_clk;
  assign mem_190_5_R0_en = R0_en & R0_addr_sel == 8'hbe;
  assign mem_190_5_W0_addr = W0_addr[25:0];
  assign mem_190_5_W0_clk = W0_clk;
  assign mem_190_5_W0_data = W0_data[47:40];
  assign mem_190_5_W0_en = W0_en & W0_addr_sel == 8'hbe;
  assign mem_190_5_W0_mask = W0_mask[5];
  assign mem_190_6_R0_addr = R0_addr[25:0];
  assign mem_190_6_R0_clk = R0_clk;
  assign mem_190_6_R0_en = R0_en & R0_addr_sel == 8'hbe;
  assign mem_190_6_W0_addr = W0_addr[25:0];
  assign mem_190_6_W0_clk = W0_clk;
  assign mem_190_6_W0_data = W0_data[55:48];
  assign mem_190_6_W0_en = W0_en & W0_addr_sel == 8'hbe;
  assign mem_190_6_W0_mask = W0_mask[6];
  assign mem_190_7_R0_addr = R0_addr[25:0];
  assign mem_190_7_R0_clk = R0_clk;
  assign mem_190_7_R0_en = R0_en & R0_addr_sel == 8'hbe;
  assign mem_190_7_W0_addr = W0_addr[25:0];
  assign mem_190_7_W0_clk = W0_clk;
  assign mem_190_7_W0_data = W0_data[63:56];
  assign mem_190_7_W0_en = W0_en & W0_addr_sel == 8'hbe;
  assign mem_190_7_W0_mask = W0_mask[7];
  assign mem_191_0_R0_addr = R0_addr[25:0];
  assign mem_191_0_R0_clk = R0_clk;
  assign mem_191_0_R0_en = R0_en & R0_addr_sel == 8'hbf;
  assign mem_191_0_W0_addr = W0_addr[25:0];
  assign mem_191_0_W0_clk = W0_clk;
  assign mem_191_0_W0_data = W0_data[7:0];
  assign mem_191_0_W0_en = W0_en & W0_addr_sel == 8'hbf;
  assign mem_191_0_W0_mask = W0_mask[0];
  assign mem_191_1_R0_addr = R0_addr[25:0];
  assign mem_191_1_R0_clk = R0_clk;
  assign mem_191_1_R0_en = R0_en & R0_addr_sel == 8'hbf;
  assign mem_191_1_W0_addr = W0_addr[25:0];
  assign mem_191_1_W0_clk = W0_clk;
  assign mem_191_1_W0_data = W0_data[15:8];
  assign mem_191_1_W0_en = W0_en & W0_addr_sel == 8'hbf;
  assign mem_191_1_W0_mask = W0_mask[1];
  assign mem_191_2_R0_addr = R0_addr[25:0];
  assign mem_191_2_R0_clk = R0_clk;
  assign mem_191_2_R0_en = R0_en & R0_addr_sel == 8'hbf;
  assign mem_191_2_W0_addr = W0_addr[25:0];
  assign mem_191_2_W0_clk = W0_clk;
  assign mem_191_2_W0_data = W0_data[23:16];
  assign mem_191_2_W0_en = W0_en & W0_addr_sel == 8'hbf;
  assign mem_191_2_W0_mask = W0_mask[2];
  assign mem_191_3_R0_addr = R0_addr[25:0];
  assign mem_191_3_R0_clk = R0_clk;
  assign mem_191_3_R0_en = R0_en & R0_addr_sel == 8'hbf;
  assign mem_191_3_W0_addr = W0_addr[25:0];
  assign mem_191_3_W0_clk = W0_clk;
  assign mem_191_3_W0_data = W0_data[31:24];
  assign mem_191_3_W0_en = W0_en & W0_addr_sel == 8'hbf;
  assign mem_191_3_W0_mask = W0_mask[3];
  assign mem_191_4_R0_addr = R0_addr[25:0];
  assign mem_191_4_R0_clk = R0_clk;
  assign mem_191_4_R0_en = R0_en & R0_addr_sel == 8'hbf;
  assign mem_191_4_W0_addr = W0_addr[25:0];
  assign mem_191_4_W0_clk = W0_clk;
  assign mem_191_4_W0_data = W0_data[39:32];
  assign mem_191_4_W0_en = W0_en & W0_addr_sel == 8'hbf;
  assign mem_191_4_W0_mask = W0_mask[4];
  assign mem_191_5_R0_addr = R0_addr[25:0];
  assign mem_191_5_R0_clk = R0_clk;
  assign mem_191_5_R0_en = R0_en & R0_addr_sel == 8'hbf;
  assign mem_191_5_W0_addr = W0_addr[25:0];
  assign mem_191_5_W0_clk = W0_clk;
  assign mem_191_5_W0_data = W0_data[47:40];
  assign mem_191_5_W0_en = W0_en & W0_addr_sel == 8'hbf;
  assign mem_191_5_W0_mask = W0_mask[5];
  assign mem_191_6_R0_addr = R0_addr[25:0];
  assign mem_191_6_R0_clk = R0_clk;
  assign mem_191_6_R0_en = R0_en & R0_addr_sel == 8'hbf;
  assign mem_191_6_W0_addr = W0_addr[25:0];
  assign mem_191_6_W0_clk = W0_clk;
  assign mem_191_6_W0_data = W0_data[55:48];
  assign mem_191_6_W0_en = W0_en & W0_addr_sel == 8'hbf;
  assign mem_191_6_W0_mask = W0_mask[6];
  assign mem_191_7_R0_addr = R0_addr[25:0];
  assign mem_191_7_R0_clk = R0_clk;
  assign mem_191_7_R0_en = R0_en & R0_addr_sel == 8'hbf;
  assign mem_191_7_W0_addr = W0_addr[25:0];
  assign mem_191_7_W0_clk = W0_clk;
  assign mem_191_7_W0_data = W0_data[63:56];
  assign mem_191_7_W0_en = W0_en & W0_addr_sel == 8'hbf;
  assign mem_191_7_W0_mask = W0_mask[7];
  assign mem_192_0_R0_addr = R0_addr[25:0];
  assign mem_192_0_R0_clk = R0_clk;
  assign mem_192_0_R0_en = R0_en & R0_addr_sel == 8'hc0;
  assign mem_192_0_W0_addr = W0_addr[25:0];
  assign mem_192_0_W0_clk = W0_clk;
  assign mem_192_0_W0_data = W0_data[7:0];
  assign mem_192_0_W0_en = W0_en & W0_addr_sel == 8'hc0;
  assign mem_192_0_W0_mask = W0_mask[0];
  assign mem_192_1_R0_addr = R0_addr[25:0];
  assign mem_192_1_R0_clk = R0_clk;
  assign mem_192_1_R0_en = R0_en & R0_addr_sel == 8'hc0;
  assign mem_192_1_W0_addr = W0_addr[25:0];
  assign mem_192_1_W0_clk = W0_clk;
  assign mem_192_1_W0_data = W0_data[15:8];
  assign mem_192_1_W0_en = W0_en & W0_addr_sel == 8'hc0;
  assign mem_192_1_W0_mask = W0_mask[1];
  assign mem_192_2_R0_addr = R0_addr[25:0];
  assign mem_192_2_R0_clk = R0_clk;
  assign mem_192_2_R0_en = R0_en & R0_addr_sel == 8'hc0;
  assign mem_192_2_W0_addr = W0_addr[25:0];
  assign mem_192_2_W0_clk = W0_clk;
  assign mem_192_2_W0_data = W0_data[23:16];
  assign mem_192_2_W0_en = W0_en & W0_addr_sel == 8'hc0;
  assign mem_192_2_W0_mask = W0_mask[2];
  assign mem_192_3_R0_addr = R0_addr[25:0];
  assign mem_192_3_R0_clk = R0_clk;
  assign mem_192_3_R0_en = R0_en & R0_addr_sel == 8'hc0;
  assign mem_192_3_W0_addr = W0_addr[25:0];
  assign mem_192_3_W0_clk = W0_clk;
  assign mem_192_3_W0_data = W0_data[31:24];
  assign mem_192_3_W0_en = W0_en & W0_addr_sel == 8'hc0;
  assign mem_192_3_W0_mask = W0_mask[3];
  assign mem_192_4_R0_addr = R0_addr[25:0];
  assign mem_192_4_R0_clk = R0_clk;
  assign mem_192_4_R0_en = R0_en & R0_addr_sel == 8'hc0;
  assign mem_192_4_W0_addr = W0_addr[25:0];
  assign mem_192_4_W0_clk = W0_clk;
  assign mem_192_4_W0_data = W0_data[39:32];
  assign mem_192_4_W0_en = W0_en & W0_addr_sel == 8'hc0;
  assign mem_192_4_W0_mask = W0_mask[4];
  assign mem_192_5_R0_addr = R0_addr[25:0];
  assign mem_192_5_R0_clk = R0_clk;
  assign mem_192_5_R0_en = R0_en & R0_addr_sel == 8'hc0;
  assign mem_192_5_W0_addr = W0_addr[25:0];
  assign mem_192_5_W0_clk = W0_clk;
  assign mem_192_5_W0_data = W0_data[47:40];
  assign mem_192_5_W0_en = W0_en & W0_addr_sel == 8'hc0;
  assign mem_192_5_W0_mask = W0_mask[5];
  assign mem_192_6_R0_addr = R0_addr[25:0];
  assign mem_192_6_R0_clk = R0_clk;
  assign mem_192_6_R0_en = R0_en & R0_addr_sel == 8'hc0;
  assign mem_192_6_W0_addr = W0_addr[25:0];
  assign mem_192_6_W0_clk = W0_clk;
  assign mem_192_6_W0_data = W0_data[55:48];
  assign mem_192_6_W0_en = W0_en & W0_addr_sel == 8'hc0;
  assign mem_192_6_W0_mask = W0_mask[6];
  assign mem_192_7_R0_addr = R0_addr[25:0];
  assign mem_192_7_R0_clk = R0_clk;
  assign mem_192_7_R0_en = R0_en & R0_addr_sel == 8'hc0;
  assign mem_192_7_W0_addr = W0_addr[25:0];
  assign mem_192_7_W0_clk = W0_clk;
  assign mem_192_7_W0_data = W0_data[63:56];
  assign mem_192_7_W0_en = W0_en & W0_addr_sel == 8'hc0;
  assign mem_192_7_W0_mask = W0_mask[7];
  assign mem_193_0_R0_addr = R0_addr[25:0];
  assign mem_193_0_R0_clk = R0_clk;
  assign mem_193_0_R0_en = R0_en & R0_addr_sel == 8'hc1;
  assign mem_193_0_W0_addr = W0_addr[25:0];
  assign mem_193_0_W0_clk = W0_clk;
  assign mem_193_0_W0_data = W0_data[7:0];
  assign mem_193_0_W0_en = W0_en & W0_addr_sel == 8'hc1;
  assign mem_193_0_W0_mask = W0_mask[0];
  assign mem_193_1_R0_addr = R0_addr[25:0];
  assign mem_193_1_R0_clk = R0_clk;
  assign mem_193_1_R0_en = R0_en & R0_addr_sel == 8'hc1;
  assign mem_193_1_W0_addr = W0_addr[25:0];
  assign mem_193_1_W0_clk = W0_clk;
  assign mem_193_1_W0_data = W0_data[15:8];
  assign mem_193_1_W0_en = W0_en & W0_addr_sel == 8'hc1;
  assign mem_193_1_W0_mask = W0_mask[1];
  assign mem_193_2_R0_addr = R0_addr[25:0];
  assign mem_193_2_R0_clk = R0_clk;
  assign mem_193_2_R0_en = R0_en & R0_addr_sel == 8'hc1;
  assign mem_193_2_W0_addr = W0_addr[25:0];
  assign mem_193_2_W0_clk = W0_clk;
  assign mem_193_2_W0_data = W0_data[23:16];
  assign mem_193_2_W0_en = W0_en & W0_addr_sel == 8'hc1;
  assign mem_193_2_W0_mask = W0_mask[2];
  assign mem_193_3_R0_addr = R0_addr[25:0];
  assign mem_193_3_R0_clk = R0_clk;
  assign mem_193_3_R0_en = R0_en & R0_addr_sel == 8'hc1;
  assign mem_193_3_W0_addr = W0_addr[25:0];
  assign mem_193_3_W0_clk = W0_clk;
  assign mem_193_3_W0_data = W0_data[31:24];
  assign mem_193_3_W0_en = W0_en & W0_addr_sel == 8'hc1;
  assign mem_193_3_W0_mask = W0_mask[3];
  assign mem_193_4_R0_addr = R0_addr[25:0];
  assign mem_193_4_R0_clk = R0_clk;
  assign mem_193_4_R0_en = R0_en & R0_addr_sel == 8'hc1;
  assign mem_193_4_W0_addr = W0_addr[25:0];
  assign mem_193_4_W0_clk = W0_clk;
  assign mem_193_4_W0_data = W0_data[39:32];
  assign mem_193_4_W0_en = W0_en & W0_addr_sel == 8'hc1;
  assign mem_193_4_W0_mask = W0_mask[4];
  assign mem_193_5_R0_addr = R0_addr[25:0];
  assign mem_193_5_R0_clk = R0_clk;
  assign mem_193_5_R0_en = R0_en & R0_addr_sel == 8'hc1;
  assign mem_193_5_W0_addr = W0_addr[25:0];
  assign mem_193_5_W0_clk = W0_clk;
  assign mem_193_5_W0_data = W0_data[47:40];
  assign mem_193_5_W0_en = W0_en & W0_addr_sel == 8'hc1;
  assign mem_193_5_W0_mask = W0_mask[5];
  assign mem_193_6_R0_addr = R0_addr[25:0];
  assign mem_193_6_R0_clk = R0_clk;
  assign mem_193_6_R0_en = R0_en & R0_addr_sel == 8'hc1;
  assign mem_193_6_W0_addr = W0_addr[25:0];
  assign mem_193_6_W0_clk = W0_clk;
  assign mem_193_6_W0_data = W0_data[55:48];
  assign mem_193_6_W0_en = W0_en & W0_addr_sel == 8'hc1;
  assign mem_193_6_W0_mask = W0_mask[6];
  assign mem_193_7_R0_addr = R0_addr[25:0];
  assign mem_193_7_R0_clk = R0_clk;
  assign mem_193_7_R0_en = R0_en & R0_addr_sel == 8'hc1;
  assign mem_193_7_W0_addr = W0_addr[25:0];
  assign mem_193_7_W0_clk = W0_clk;
  assign mem_193_7_W0_data = W0_data[63:56];
  assign mem_193_7_W0_en = W0_en & W0_addr_sel == 8'hc1;
  assign mem_193_7_W0_mask = W0_mask[7];
  assign mem_194_0_R0_addr = R0_addr[25:0];
  assign mem_194_0_R0_clk = R0_clk;
  assign mem_194_0_R0_en = R0_en & R0_addr_sel == 8'hc2;
  assign mem_194_0_W0_addr = W0_addr[25:0];
  assign mem_194_0_W0_clk = W0_clk;
  assign mem_194_0_W0_data = W0_data[7:0];
  assign mem_194_0_W0_en = W0_en & W0_addr_sel == 8'hc2;
  assign mem_194_0_W0_mask = W0_mask[0];
  assign mem_194_1_R0_addr = R0_addr[25:0];
  assign mem_194_1_R0_clk = R0_clk;
  assign mem_194_1_R0_en = R0_en & R0_addr_sel == 8'hc2;
  assign mem_194_1_W0_addr = W0_addr[25:0];
  assign mem_194_1_W0_clk = W0_clk;
  assign mem_194_1_W0_data = W0_data[15:8];
  assign mem_194_1_W0_en = W0_en & W0_addr_sel == 8'hc2;
  assign mem_194_1_W0_mask = W0_mask[1];
  assign mem_194_2_R0_addr = R0_addr[25:0];
  assign mem_194_2_R0_clk = R0_clk;
  assign mem_194_2_R0_en = R0_en & R0_addr_sel == 8'hc2;
  assign mem_194_2_W0_addr = W0_addr[25:0];
  assign mem_194_2_W0_clk = W0_clk;
  assign mem_194_2_W0_data = W0_data[23:16];
  assign mem_194_2_W0_en = W0_en & W0_addr_sel == 8'hc2;
  assign mem_194_2_W0_mask = W0_mask[2];
  assign mem_194_3_R0_addr = R0_addr[25:0];
  assign mem_194_3_R0_clk = R0_clk;
  assign mem_194_3_R0_en = R0_en & R0_addr_sel == 8'hc2;
  assign mem_194_3_W0_addr = W0_addr[25:0];
  assign mem_194_3_W0_clk = W0_clk;
  assign mem_194_3_W0_data = W0_data[31:24];
  assign mem_194_3_W0_en = W0_en & W0_addr_sel == 8'hc2;
  assign mem_194_3_W0_mask = W0_mask[3];
  assign mem_194_4_R0_addr = R0_addr[25:0];
  assign mem_194_4_R0_clk = R0_clk;
  assign mem_194_4_R0_en = R0_en & R0_addr_sel == 8'hc2;
  assign mem_194_4_W0_addr = W0_addr[25:0];
  assign mem_194_4_W0_clk = W0_clk;
  assign mem_194_4_W0_data = W0_data[39:32];
  assign mem_194_4_W0_en = W0_en & W0_addr_sel == 8'hc2;
  assign mem_194_4_W0_mask = W0_mask[4];
  assign mem_194_5_R0_addr = R0_addr[25:0];
  assign mem_194_5_R0_clk = R0_clk;
  assign mem_194_5_R0_en = R0_en & R0_addr_sel == 8'hc2;
  assign mem_194_5_W0_addr = W0_addr[25:0];
  assign mem_194_5_W0_clk = W0_clk;
  assign mem_194_5_W0_data = W0_data[47:40];
  assign mem_194_5_W0_en = W0_en & W0_addr_sel == 8'hc2;
  assign mem_194_5_W0_mask = W0_mask[5];
  assign mem_194_6_R0_addr = R0_addr[25:0];
  assign mem_194_6_R0_clk = R0_clk;
  assign mem_194_6_R0_en = R0_en & R0_addr_sel == 8'hc2;
  assign mem_194_6_W0_addr = W0_addr[25:0];
  assign mem_194_6_W0_clk = W0_clk;
  assign mem_194_6_W0_data = W0_data[55:48];
  assign mem_194_6_W0_en = W0_en & W0_addr_sel == 8'hc2;
  assign mem_194_6_W0_mask = W0_mask[6];
  assign mem_194_7_R0_addr = R0_addr[25:0];
  assign mem_194_7_R0_clk = R0_clk;
  assign mem_194_7_R0_en = R0_en & R0_addr_sel == 8'hc2;
  assign mem_194_7_W0_addr = W0_addr[25:0];
  assign mem_194_7_W0_clk = W0_clk;
  assign mem_194_7_W0_data = W0_data[63:56];
  assign mem_194_7_W0_en = W0_en & W0_addr_sel == 8'hc2;
  assign mem_194_7_W0_mask = W0_mask[7];
  assign mem_195_0_R0_addr = R0_addr[25:0];
  assign mem_195_0_R0_clk = R0_clk;
  assign mem_195_0_R0_en = R0_en & R0_addr_sel == 8'hc3;
  assign mem_195_0_W0_addr = W0_addr[25:0];
  assign mem_195_0_W0_clk = W0_clk;
  assign mem_195_0_W0_data = W0_data[7:0];
  assign mem_195_0_W0_en = W0_en & W0_addr_sel == 8'hc3;
  assign mem_195_0_W0_mask = W0_mask[0];
  assign mem_195_1_R0_addr = R0_addr[25:0];
  assign mem_195_1_R0_clk = R0_clk;
  assign mem_195_1_R0_en = R0_en & R0_addr_sel == 8'hc3;
  assign mem_195_1_W0_addr = W0_addr[25:0];
  assign mem_195_1_W0_clk = W0_clk;
  assign mem_195_1_W0_data = W0_data[15:8];
  assign mem_195_1_W0_en = W0_en & W0_addr_sel == 8'hc3;
  assign mem_195_1_W0_mask = W0_mask[1];
  assign mem_195_2_R0_addr = R0_addr[25:0];
  assign mem_195_2_R0_clk = R0_clk;
  assign mem_195_2_R0_en = R0_en & R0_addr_sel == 8'hc3;
  assign mem_195_2_W0_addr = W0_addr[25:0];
  assign mem_195_2_W0_clk = W0_clk;
  assign mem_195_2_W0_data = W0_data[23:16];
  assign mem_195_2_W0_en = W0_en & W0_addr_sel == 8'hc3;
  assign mem_195_2_W0_mask = W0_mask[2];
  assign mem_195_3_R0_addr = R0_addr[25:0];
  assign mem_195_3_R0_clk = R0_clk;
  assign mem_195_3_R0_en = R0_en & R0_addr_sel == 8'hc3;
  assign mem_195_3_W0_addr = W0_addr[25:0];
  assign mem_195_3_W0_clk = W0_clk;
  assign mem_195_3_W0_data = W0_data[31:24];
  assign mem_195_3_W0_en = W0_en & W0_addr_sel == 8'hc3;
  assign mem_195_3_W0_mask = W0_mask[3];
  assign mem_195_4_R0_addr = R0_addr[25:0];
  assign mem_195_4_R0_clk = R0_clk;
  assign mem_195_4_R0_en = R0_en & R0_addr_sel == 8'hc3;
  assign mem_195_4_W0_addr = W0_addr[25:0];
  assign mem_195_4_W0_clk = W0_clk;
  assign mem_195_4_W0_data = W0_data[39:32];
  assign mem_195_4_W0_en = W0_en & W0_addr_sel == 8'hc3;
  assign mem_195_4_W0_mask = W0_mask[4];
  assign mem_195_5_R0_addr = R0_addr[25:0];
  assign mem_195_5_R0_clk = R0_clk;
  assign mem_195_5_R0_en = R0_en & R0_addr_sel == 8'hc3;
  assign mem_195_5_W0_addr = W0_addr[25:0];
  assign mem_195_5_W0_clk = W0_clk;
  assign mem_195_5_W0_data = W0_data[47:40];
  assign mem_195_5_W0_en = W0_en & W0_addr_sel == 8'hc3;
  assign mem_195_5_W0_mask = W0_mask[5];
  assign mem_195_6_R0_addr = R0_addr[25:0];
  assign mem_195_6_R0_clk = R0_clk;
  assign mem_195_6_R0_en = R0_en & R0_addr_sel == 8'hc3;
  assign mem_195_6_W0_addr = W0_addr[25:0];
  assign mem_195_6_W0_clk = W0_clk;
  assign mem_195_6_W0_data = W0_data[55:48];
  assign mem_195_6_W0_en = W0_en & W0_addr_sel == 8'hc3;
  assign mem_195_6_W0_mask = W0_mask[6];
  assign mem_195_7_R0_addr = R0_addr[25:0];
  assign mem_195_7_R0_clk = R0_clk;
  assign mem_195_7_R0_en = R0_en & R0_addr_sel == 8'hc3;
  assign mem_195_7_W0_addr = W0_addr[25:0];
  assign mem_195_7_W0_clk = W0_clk;
  assign mem_195_7_W0_data = W0_data[63:56];
  assign mem_195_7_W0_en = W0_en & W0_addr_sel == 8'hc3;
  assign mem_195_7_W0_mask = W0_mask[7];
  assign mem_196_0_R0_addr = R0_addr[25:0];
  assign mem_196_0_R0_clk = R0_clk;
  assign mem_196_0_R0_en = R0_en & R0_addr_sel == 8'hc4;
  assign mem_196_0_W0_addr = W0_addr[25:0];
  assign mem_196_0_W0_clk = W0_clk;
  assign mem_196_0_W0_data = W0_data[7:0];
  assign mem_196_0_W0_en = W0_en & W0_addr_sel == 8'hc4;
  assign mem_196_0_W0_mask = W0_mask[0];
  assign mem_196_1_R0_addr = R0_addr[25:0];
  assign mem_196_1_R0_clk = R0_clk;
  assign mem_196_1_R0_en = R0_en & R0_addr_sel == 8'hc4;
  assign mem_196_1_W0_addr = W0_addr[25:0];
  assign mem_196_1_W0_clk = W0_clk;
  assign mem_196_1_W0_data = W0_data[15:8];
  assign mem_196_1_W0_en = W0_en & W0_addr_sel == 8'hc4;
  assign mem_196_1_W0_mask = W0_mask[1];
  assign mem_196_2_R0_addr = R0_addr[25:0];
  assign mem_196_2_R0_clk = R0_clk;
  assign mem_196_2_R0_en = R0_en & R0_addr_sel == 8'hc4;
  assign mem_196_2_W0_addr = W0_addr[25:0];
  assign mem_196_2_W0_clk = W0_clk;
  assign mem_196_2_W0_data = W0_data[23:16];
  assign mem_196_2_W0_en = W0_en & W0_addr_sel == 8'hc4;
  assign mem_196_2_W0_mask = W0_mask[2];
  assign mem_196_3_R0_addr = R0_addr[25:0];
  assign mem_196_3_R0_clk = R0_clk;
  assign mem_196_3_R0_en = R0_en & R0_addr_sel == 8'hc4;
  assign mem_196_3_W0_addr = W0_addr[25:0];
  assign mem_196_3_W0_clk = W0_clk;
  assign mem_196_3_W0_data = W0_data[31:24];
  assign mem_196_3_W0_en = W0_en & W0_addr_sel == 8'hc4;
  assign mem_196_3_W0_mask = W0_mask[3];
  assign mem_196_4_R0_addr = R0_addr[25:0];
  assign mem_196_4_R0_clk = R0_clk;
  assign mem_196_4_R0_en = R0_en & R0_addr_sel == 8'hc4;
  assign mem_196_4_W0_addr = W0_addr[25:0];
  assign mem_196_4_W0_clk = W0_clk;
  assign mem_196_4_W0_data = W0_data[39:32];
  assign mem_196_4_W0_en = W0_en & W0_addr_sel == 8'hc4;
  assign mem_196_4_W0_mask = W0_mask[4];
  assign mem_196_5_R0_addr = R0_addr[25:0];
  assign mem_196_5_R0_clk = R0_clk;
  assign mem_196_5_R0_en = R0_en & R0_addr_sel == 8'hc4;
  assign mem_196_5_W0_addr = W0_addr[25:0];
  assign mem_196_5_W0_clk = W0_clk;
  assign mem_196_5_W0_data = W0_data[47:40];
  assign mem_196_5_W0_en = W0_en & W0_addr_sel == 8'hc4;
  assign mem_196_5_W0_mask = W0_mask[5];
  assign mem_196_6_R0_addr = R0_addr[25:0];
  assign mem_196_6_R0_clk = R0_clk;
  assign mem_196_6_R0_en = R0_en & R0_addr_sel == 8'hc4;
  assign mem_196_6_W0_addr = W0_addr[25:0];
  assign mem_196_6_W0_clk = W0_clk;
  assign mem_196_6_W0_data = W0_data[55:48];
  assign mem_196_6_W0_en = W0_en & W0_addr_sel == 8'hc4;
  assign mem_196_6_W0_mask = W0_mask[6];
  assign mem_196_7_R0_addr = R0_addr[25:0];
  assign mem_196_7_R0_clk = R0_clk;
  assign mem_196_7_R0_en = R0_en & R0_addr_sel == 8'hc4;
  assign mem_196_7_W0_addr = W0_addr[25:0];
  assign mem_196_7_W0_clk = W0_clk;
  assign mem_196_7_W0_data = W0_data[63:56];
  assign mem_196_7_W0_en = W0_en & W0_addr_sel == 8'hc4;
  assign mem_196_7_W0_mask = W0_mask[7];
  assign mem_197_0_R0_addr = R0_addr[25:0];
  assign mem_197_0_R0_clk = R0_clk;
  assign mem_197_0_R0_en = R0_en & R0_addr_sel == 8'hc5;
  assign mem_197_0_W0_addr = W0_addr[25:0];
  assign mem_197_0_W0_clk = W0_clk;
  assign mem_197_0_W0_data = W0_data[7:0];
  assign mem_197_0_W0_en = W0_en & W0_addr_sel == 8'hc5;
  assign mem_197_0_W0_mask = W0_mask[0];
  assign mem_197_1_R0_addr = R0_addr[25:0];
  assign mem_197_1_R0_clk = R0_clk;
  assign mem_197_1_R0_en = R0_en & R0_addr_sel == 8'hc5;
  assign mem_197_1_W0_addr = W0_addr[25:0];
  assign mem_197_1_W0_clk = W0_clk;
  assign mem_197_1_W0_data = W0_data[15:8];
  assign mem_197_1_W0_en = W0_en & W0_addr_sel == 8'hc5;
  assign mem_197_1_W0_mask = W0_mask[1];
  assign mem_197_2_R0_addr = R0_addr[25:0];
  assign mem_197_2_R0_clk = R0_clk;
  assign mem_197_2_R0_en = R0_en & R0_addr_sel == 8'hc5;
  assign mem_197_2_W0_addr = W0_addr[25:0];
  assign mem_197_2_W0_clk = W0_clk;
  assign mem_197_2_W0_data = W0_data[23:16];
  assign mem_197_2_W0_en = W0_en & W0_addr_sel == 8'hc5;
  assign mem_197_2_W0_mask = W0_mask[2];
  assign mem_197_3_R0_addr = R0_addr[25:0];
  assign mem_197_3_R0_clk = R0_clk;
  assign mem_197_3_R0_en = R0_en & R0_addr_sel == 8'hc5;
  assign mem_197_3_W0_addr = W0_addr[25:0];
  assign mem_197_3_W0_clk = W0_clk;
  assign mem_197_3_W0_data = W0_data[31:24];
  assign mem_197_3_W0_en = W0_en & W0_addr_sel == 8'hc5;
  assign mem_197_3_W0_mask = W0_mask[3];
  assign mem_197_4_R0_addr = R0_addr[25:0];
  assign mem_197_4_R0_clk = R0_clk;
  assign mem_197_4_R0_en = R0_en & R0_addr_sel == 8'hc5;
  assign mem_197_4_W0_addr = W0_addr[25:0];
  assign mem_197_4_W0_clk = W0_clk;
  assign mem_197_4_W0_data = W0_data[39:32];
  assign mem_197_4_W0_en = W0_en & W0_addr_sel == 8'hc5;
  assign mem_197_4_W0_mask = W0_mask[4];
  assign mem_197_5_R0_addr = R0_addr[25:0];
  assign mem_197_5_R0_clk = R0_clk;
  assign mem_197_5_R0_en = R0_en & R0_addr_sel == 8'hc5;
  assign mem_197_5_W0_addr = W0_addr[25:0];
  assign mem_197_5_W0_clk = W0_clk;
  assign mem_197_5_W0_data = W0_data[47:40];
  assign mem_197_5_W0_en = W0_en & W0_addr_sel == 8'hc5;
  assign mem_197_5_W0_mask = W0_mask[5];
  assign mem_197_6_R0_addr = R0_addr[25:0];
  assign mem_197_6_R0_clk = R0_clk;
  assign mem_197_6_R0_en = R0_en & R0_addr_sel == 8'hc5;
  assign mem_197_6_W0_addr = W0_addr[25:0];
  assign mem_197_6_W0_clk = W0_clk;
  assign mem_197_6_W0_data = W0_data[55:48];
  assign mem_197_6_W0_en = W0_en & W0_addr_sel == 8'hc5;
  assign mem_197_6_W0_mask = W0_mask[6];
  assign mem_197_7_R0_addr = R0_addr[25:0];
  assign mem_197_7_R0_clk = R0_clk;
  assign mem_197_7_R0_en = R0_en & R0_addr_sel == 8'hc5;
  assign mem_197_7_W0_addr = W0_addr[25:0];
  assign mem_197_7_W0_clk = W0_clk;
  assign mem_197_7_W0_data = W0_data[63:56];
  assign mem_197_7_W0_en = W0_en & W0_addr_sel == 8'hc5;
  assign mem_197_7_W0_mask = W0_mask[7];
  assign mem_198_0_R0_addr = R0_addr[25:0];
  assign mem_198_0_R0_clk = R0_clk;
  assign mem_198_0_R0_en = R0_en & R0_addr_sel == 8'hc6;
  assign mem_198_0_W0_addr = W0_addr[25:0];
  assign mem_198_0_W0_clk = W0_clk;
  assign mem_198_0_W0_data = W0_data[7:0];
  assign mem_198_0_W0_en = W0_en & W0_addr_sel == 8'hc6;
  assign mem_198_0_W0_mask = W0_mask[0];
  assign mem_198_1_R0_addr = R0_addr[25:0];
  assign mem_198_1_R0_clk = R0_clk;
  assign mem_198_1_R0_en = R0_en & R0_addr_sel == 8'hc6;
  assign mem_198_1_W0_addr = W0_addr[25:0];
  assign mem_198_1_W0_clk = W0_clk;
  assign mem_198_1_W0_data = W0_data[15:8];
  assign mem_198_1_W0_en = W0_en & W0_addr_sel == 8'hc6;
  assign mem_198_1_W0_mask = W0_mask[1];
  assign mem_198_2_R0_addr = R0_addr[25:0];
  assign mem_198_2_R0_clk = R0_clk;
  assign mem_198_2_R0_en = R0_en & R0_addr_sel == 8'hc6;
  assign mem_198_2_W0_addr = W0_addr[25:0];
  assign mem_198_2_W0_clk = W0_clk;
  assign mem_198_2_W0_data = W0_data[23:16];
  assign mem_198_2_W0_en = W0_en & W0_addr_sel == 8'hc6;
  assign mem_198_2_W0_mask = W0_mask[2];
  assign mem_198_3_R0_addr = R0_addr[25:0];
  assign mem_198_3_R0_clk = R0_clk;
  assign mem_198_3_R0_en = R0_en & R0_addr_sel == 8'hc6;
  assign mem_198_3_W0_addr = W0_addr[25:0];
  assign mem_198_3_W0_clk = W0_clk;
  assign mem_198_3_W0_data = W0_data[31:24];
  assign mem_198_3_W0_en = W0_en & W0_addr_sel == 8'hc6;
  assign mem_198_3_W0_mask = W0_mask[3];
  assign mem_198_4_R0_addr = R0_addr[25:0];
  assign mem_198_4_R0_clk = R0_clk;
  assign mem_198_4_R0_en = R0_en & R0_addr_sel == 8'hc6;
  assign mem_198_4_W0_addr = W0_addr[25:0];
  assign mem_198_4_W0_clk = W0_clk;
  assign mem_198_4_W0_data = W0_data[39:32];
  assign mem_198_4_W0_en = W0_en & W0_addr_sel == 8'hc6;
  assign mem_198_4_W0_mask = W0_mask[4];
  assign mem_198_5_R0_addr = R0_addr[25:0];
  assign mem_198_5_R0_clk = R0_clk;
  assign mem_198_5_R0_en = R0_en & R0_addr_sel == 8'hc6;
  assign mem_198_5_W0_addr = W0_addr[25:0];
  assign mem_198_5_W0_clk = W0_clk;
  assign mem_198_5_W0_data = W0_data[47:40];
  assign mem_198_5_W0_en = W0_en & W0_addr_sel == 8'hc6;
  assign mem_198_5_W0_mask = W0_mask[5];
  assign mem_198_6_R0_addr = R0_addr[25:0];
  assign mem_198_6_R0_clk = R0_clk;
  assign mem_198_6_R0_en = R0_en & R0_addr_sel == 8'hc6;
  assign mem_198_6_W0_addr = W0_addr[25:0];
  assign mem_198_6_W0_clk = W0_clk;
  assign mem_198_6_W0_data = W0_data[55:48];
  assign mem_198_6_W0_en = W0_en & W0_addr_sel == 8'hc6;
  assign mem_198_6_W0_mask = W0_mask[6];
  assign mem_198_7_R0_addr = R0_addr[25:0];
  assign mem_198_7_R0_clk = R0_clk;
  assign mem_198_7_R0_en = R0_en & R0_addr_sel == 8'hc6;
  assign mem_198_7_W0_addr = W0_addr[25:0];
  assign mem_198_7_W0_clk = W0_clk;
  assign mem_198_7_W0_data = W0_data[63:56];
  assign mem_198_7_W0_en = W0_en & W0_addr_sel == 8'hc6;
  assign mem_198_7_W0_mask = W0_mask[7];
  assign mem_199_0_R0_addr = R0_addr[25:0];
  assign mem_199_0_R0_clk = R0_clk;
  assign mem_199_0_R0_en = R0_en & R0_addr_sel == 8'hc7;
  assign mem_199_0_W0_addr = W0_addr[25:0];
  assign mem_199_0_W0_clk = W0_clk;
  assign mem_199_0_W0_data = W0_data[7:0];
  assign mem_199_0_W0_en = W0_en & W0_addr_sel == 8'hc7;
  assign mem_199_0_W0_mask = W0_mask[0];
  assign mem_199_1_R0_addr = R0_addr[25:0];
  assign mem_199_1_R0_clk = R0_clk;
  assign mem_199_1_R0_en = R0_en & R0_addr_sel == 8'hc7;
  assign mem_199_1_W0_addr = W0_addr[25:0];
  assign mem_199_1_W0_clk = W0_clk;
  assign mem_199_1_W0_data = W0_data[15:8];
  assign mem_199_1_W0_en = W0_en & W0_addr_sel == 8'hc7;
  assign mem_199_1_W0_mask = W0_mask[1];
  assign mem_199_2_R0_addr = R0_addr[25:0];
  assign mem_199_2_R0_clk = R0_clk;
  assign mem_199_2_R0_en = R0_en & R0_addr_sel == 8'hc7;
  assign mem_199_2_W0_addr = W0_addr[25:0];
  assign mem_199_2_W0_clk = W0_clk;
  assign mem_199_2_W0_data = W0_data[23:16];
  assign mem_199_2_W0_en = W0_en & W0_addr_sel == 8'hc7;
  assign mem_199_2_W0_mask = W0_mask[2];
  assign mem_199_3_R0_addr = R0_addr[25:0];
  assign mem_199_3_R0_clk = R0_clk;
  assign mem_199_3_R0_en = R0_en & R0_addr_sel == 8'hc7;
  assign mem_199_3_W0_addr = W0_addr[25:0];
  assign mem_199_3_W0_clk = W0_clk;
  assign mem_199_3_W0_data = W0_data[31:24];
  assign mem_199_3_W0_en = W0_en & W0_addr_sel == 8'hc7;
  assign mem_199_3_W0_mask = W0_mask[3];
  assign mem_199_4_R0_addr = R0_addr[25:0];
  assign mem_199_4_R0_clk = R0_clk;
  assign mem_199_4_R0_en = R0_en & R0_addr_sel == 8'hc7;
  assign mem_199_4_W0_addr = W0_addr[25:0];
  assign mem_199_4_W0_clk = W0_clk;
  assign mem_199_4_W0_data = W0_data[39:32];
  assign mem_199_4_W0_en = W0_en & W0_addr_sel == 8'hc7;
  assign mem_199_4_W0_mask = W0_mask[4];
  assign mem_199_5_R0_addr = R0_addr[25:0];
  assign mem_199_5_R0_clk = R0_clk;
  assign mem_199_5_R0_en = R0_en & R0_addr_sel == 8'hc7;
  assign mem_199_5_W0_addr = W0_addr[25:0];
  assign mem_199_5_W0_clk = W0_clk;
  assign mem_199_5_W0_data = W0_data[47:40];
  assign mem_199_5_W0_en = W0_en & W0_addr_sel == 8'hc7;
  assign mem_199_5_W0_mask = W0_mask[5];
  assign mem_199_6_R0_addr = R0_addr[25:0];
  assign mem_199_6_R0_clk = R0_clk;
  assign mem_199_6_R0_en = R0_en & R0_addr_sel == 8'hc7;
  assign mem_199_6_W0_addr = W0_addr[25:0];
  assign mem_199_6_W0_clk = W0_clk;
  assign mem_199_6_W0_data = W0_data[55:48];
  assign mem_199_6_W0_en = W0_en & W0_addr_sel == 8'hc7;
  assign mem_199_6_W0_mask = W0_mask[6];
  assign mem_199_7_R0_addr = R0_addr[25:0];
  assign mem_199_7_R0_clk = R0_clk;
  assign mem_199_7_R0_en = R0_en & R0_addr_sel == 8'hc7;
  assign mem_199_7_W0_addr = W0_addr[25:0];
  assign mem_199_7_W0_clk = W0_clk;
  assign mem_199_7_W0_data = W0_data[63:56];
  assign mem_199_7_W0_en = W0_en & W0_addr_sel == 8'hc7;
  assign mem_199_7_W0_mask = W0_mask[7];
  assign mem_200_0_R0_addr = R0_addr[25:0];
  assign mem_200_0_R0_clk = R0_clk;
  assign mem_200_0_R0_en = R0_en & R0_addr_sel == 8'hc8;
  assign mem_200_0_W0_addr = W0_addr[25:0];
  assign mem_200_0_W0_clk = W0_clk;
  assign mem_200_0_W0_data = W0_data[7:0];
  assign mem_200_0_W0_en = W0_en & W0_addr_sel == 8'hc8;
  assign mem_200_0_W0_mask = W0_mask[0];
  assign mem_200_1_R0_addr = R0_addr[25:0];
  assign mem_200_1_R0_clk = R0_clk;
  assign mem_200_1_R0_en = R0_en & R0_addr_sel == 8'hc8;
  assign mem_200_1_W0_addr = W0_addr[25:0];
  assign mem_200_1_W0_clk = W0_clk;
  assign mem_200_1_W0_data = W0_data[15:8];
  assign mem_200_1_W0_en = W0_en & W0_addr_sel == 8'hc8;
  assign mem_200_1_W0_mask = W0_mask[1];
  assign mem_200_2_R0_addr = R0_addr[25:0];
  assign mem_200_2_R0_clk = R0_clk;
  assign mem_200_2_R0_en = R0_en & R0_addr_sel == 8'hc8;
  assign mem_200_2_W0_addr = W0_addr[25:0];
  assign mem_200_2_W0_clk = W0_clk;
  assign mem_200_2_W0_data = W0_data[23:16];
  assign mem_200_2_W0_en = W0_en & W0_addr_sel == 8'hc8;
  assign mem_200_2_W0_mask = W0_mask[2];
  assign mem_200_3_R0_addr = R0_addr[25:0];
  assign mem_200_3_R0_clk = R0_clk;
  assign mem_200_3_R0_en = R0_en & R0_addr_sel == 8'hc8;
  assign mem_200_3_W0_addr = W0_addr[25:0];
  assign mem_200_3_W0_clk = W0_clk;
  assign mem_200_3_W0_data = W0_data[31:24];
  assign mem_200_3_W0_en = W0_en & W0_addr_sel == 8'hc8;
  assign mem_200_3_W0_mask = W0_mask[3];
  assign mem_200_4_R0_addr = R0_addr[25:0];
  assign mem_200_4_R0_clk = R0_clk;
  assign mem_200_4_R0_en = R0_en & R0_addr_sel == 8'hc8;
  assign mem_200_4_W0_addr = W0_addr[25:0];
  assign mem_200_4_W0_clk = W0_clk;
  assign mem_200_4_W0_data = W0_data[39:32];
  assign mem_200_4_W0_en = W0_en & W0_addr_sel == 8'hc8;
  assign mem_200_4_W0_mask = W0_mask[4];
  assign mem_200_5_R0_addr = R0_addr[25:0];
  assign mem_200_5_R0_clk = R0_clk;
  assign mem_200_5_R0_en = R0_en & R0_addr_sel == 8'hc8;
  assign mem_200_5_W0_addr = W0_addr[25:0];
  assign mem_200_5_W0_clk = W0_clk;
  assign mem_200_5_W0_data = W0_data[47:40];
  assign mem_200_5_W0_en = W0_en & W0_addr_sel == 8'hc8;
  assign mem_200_5_W0_mask = W0_mask[5];
  assign mem_200_6_R0_addr = R0_addr[25:0];
  assign mem_200_6_R0_clk = R0_clk;
  assign mem_200_6_R0_en = R0_en & R0_addr_sel == 8'hc8;
  assign mem_200_6_W0_addr = W0_addr[25:0];
  assign mem_200_6_W0_clk = W0_clk;
  assign mem_200_6_W0_data = W0_data[55:48];
  assign mem_200_6_W0_en = W0_en & W0_addr_sel == 8'hc8;
  assign mem_200_6_W0_mask = W0_mask[6];
  assign mem_200_7_R0_addr = R0_addr[25:0];
  assign mem_200_7_R0_clk = R0_clk;
  assign mem_200_7_R0_en = R0_en & R0_addr_sel == 8'hc8;
  assign mem_200_7_W0_addr = W0_addr[25:0];
  assign mem_200_7_W0_clk = W0_clk;
  assign mem_200_7_W0_data = W0_data[63:56];
  assign mem_200_7_W0_en = W0_en & W0_addr_sel == 8'hc8;
  assign mem_200_7_W0_mask = W0_mask[7];
  assign mem_201_0_R0_addr = R0_addr[25:0];
  assign mem_201_0_R0_clk = R0_clk;
  assign mem_201_0_R0_en = R0_en & R0_addr_sel == 8'hc9;
  assign mem_201_0_W0_addr = W0_addr[25:0];
  assign mem_201_0_W0_clk = W0_clk;
  assign mem_201_0_W0_data = W0_data[7:0];
  assign mem_201_0_W0_en = W0_en & W0_addr_sel == 8'hc9;
  assign mem_201_0_W0_mask = W0_mask[0];
  assign mem_201_1_R0_addr = R0_addr[25:0];
  assign mem_201_1_R0_clk = R0_clk;
  assign mem_201_1_R0_en = R0_en & R0_addr_sel == 8'hc9;
  assign mem_201_1_W0_addr = W0_addr[25:0];
  assign mem_201_1_W0_clk = W0_clk;
  assign mem_201_1_W0_data = W0_data[15:8];
  assign mem_201_1_W0_en = W0_en & W0_addr_sel == 8'hc9;
  assign mem_201_1_W0_mask = W0_mask[1];
  assign mem_201_2_R0_addr = R0_addr[25:0];
  assign mem_201_2_R0_clk = R0_clk;
  assign mem_201_2_R0_en = R0_en & R0_addr_sel == 8'hc9;
  assign mem_201_2_W0_addr = W0_addr[25:0];
  assign mem_201_2_W0_clk = W0_clk;
  assign mem_201_2_W0_data = W0_data[23:16];
  assign mem_201_2_W0_en = W0_en & W0_addr_sel == 8'hc9;
  assign mem_201_2_W0_mask = W0_mask[2];
  assign mem_201_3_R0_addr = R0_addr[25:0];
  assign mem_201_3_R0_clk = R0_clk;
  assign mem_201_3_R0_en = R0_en & R0_addr_sel == 8'hc9;
  assign mem_201_3_W0_addr = W0_addr[25:0];
  assign mem_201_3_W0_clk = W0_clk;
  assign mem_201_3_W0_data = W0_data[31:24];
  assign mem_201_3_W0_en = W0_en & W0_addr_sel == 8'hc9;
  assign mem_201_3_W0_mask = W0_mask[3];
  assign mem_201_4_R0_addr = R0_addr[25:0];
  assign mem_201_4_R0_clk = R0_clk;
  assign mem_201_4_R0_en = R0_en & R0_addr_sel == 8'hc9;
  assign mem_201_4_W0_addr = W0_addr[25:0];
  assign mem_201_4_W0_clk = W0_clk;
  assign mem_201_4_W0_data = W0_data[39:32];
  assign mem_201_4_W0_en = W0_en & W0_addr_sel == 8'hc9;
  assign mem_201_4_W0_mask = W0_mask[4];
  assign mem_201_5_R0_addr = R0_addr[25:0];
  assign mem_201_5_R0_clk = R0_clk;
  assign mem_201_5_R0_en = R0_en & R0_addr_sel == 8'hc9;
  assign mem_201_5_W0_addr = W0_addr[25:0];
  assign mem_201_5_W0_clk = W0_clk;
  assign mem_201_5_W0_data = W0_data[47:40];
  assign mem_201_5_W0_en = W0_en & W0_addr_sel == 8'hc9;
  assign mem_201_5_W0_mask = W0_mask[5];
  assign mem_201_6_R0_addr = R0_addr[25:0];
  assign mem_201_6_R0_clk = R0_clk;
  assign mem_201_6_R0_en = R0_en & R0_addr_sel == 8'hc9;
  assign mem_201_6_W0_addr = W0_addr[25:0];
  assign mem_201_6_W0_clk = W0_clk;
  assign mem_201_6_W0_data = W0_data[55:48];
  assign mem_201_6_W0_en = W0_en & W0_addr_sel == 8'hc9;
  assign mem_201_6_W0_mask = W0_mask[6];
  assign mem_201_7_R0_addr = R0_addr[25:0];
  assign mem_201_7_R0_clk = R0_clk;
  assign mem_201_7_R0_en = R0_en & R0_addr_sel == 8'hc9;
  assign mem_201_7_W0_addr = W0_addr[25:0];
  assign mem_201_7_W0_clk = W0_clk;
  assign mem_201_7_W0_data = W0_data[63:56];
  assign mem_201_7_W0_en = W0_en & W0_addr_sel == 8'hc9;
  assign mem_201_7_W0_mask = W0_mask[7];
  assign mem_202_0_R0_addr = R0_addr[25:0];
  assign mem_202_0_R0_clk = R0_clk;
  assign mem_202_0_R0_en = R0_en & R0_addr_sel == 8'hca;
  assign mem_202_0_W0_addr = W0_addr[25:0];
  assign mem_202_0_W0_clk = W0_clk;
  assign mem_202_0_W0_data = W0_data[7:0];
  assign mem_202_0_W0_en = W0_en & W0_addr_sel == 8'hca;
  assign mem_202_0_W0_mask = W0_mask[0];
  assign mem_202_1_R0_addr = R0_addr[25:0];
  assign mem_202_1_R0_clk = R0_clk;
  assign mem_202_1_R0_en = R0_en & R0_addr_sel == 8'hca;
  assign mem_202_1_W0_addr = W0_addr[25:0];
  assign mem_202_1_W0_clk = W0_clk;
  assign mem_202_1_W0_data = W0_data[15:8];
  assign mem_202_1_W0_en = W0_en & W0_addr_sel == 8'hca;
  assign mem_202_1_W0_mask = W0_mask[1];
  assign mem_202_2_R0_addr = R0_addr[25:0];
  assign mem_202_2_R0_clk = R0_clk;
  assign mem_202_2_R0_en = R0_en & R0_addr_sel == 8'hca;
  assign mem_202_2_W0_addr = W0_addr[25:0];
  assign mem_202_2_W0_clk = W0_clk;
  assign mem_202_2_W0_data = W0_data[23:16];
  assign mem_202_2_W0_en = W0_en & W0_addr_sel == 8'hca;
  assign mem_202_2_W0_mask = W0_mask[2];
  assign mem_202_3_R0_addr = R0_addr[25:0];
  assign mem_202_3_R0_clk = R0_clk;
  assign mem_202_3_R0_en = R0_en & R0_addr_sel == 8'hca;
  assign mem_202_3_W0_addr = W0_addr[25:0];
  assign mem_202_3_W0_clk = W0_clk;
  assign mem_202_3_W0_data = W0_data[31:24];
  assign mem_202_3_W0_en = W0_en & W0_addr_sel == 8'hca;
  assign mem_202_3_W0_mask = W0_mask[3];
  assign mem_202_4_R0_addr = R0_addr[25:0];
  assign mem_202_4_R0_clk = R0_clk;
  assign mem_202_4_R0_en = R0_en & R0_addr_sel == 8'hca;
  assign mem_202_4_W0_addr = W0_addr[25:0];
  assign mem_202_4_W0_clk = W0_clk;
  assign mem_202_4_W0_data = W0_data[39:32];
  assign mem_202_4_W0_en = W0_en & W0_addr_sel == 8'hca;
  assign mem_202_4_W0_mask = W0_mask[4];
  assign mem_202_5_R0_addr = R0_addr[25:0];
  assign mem_202_5_R0_clk = R0_clk;
  assign mem_202_5_R0_en = R0_en & R0_addr_sel == 8'hca;
  assign mem_202_5_W0_addr = W0_addr[25:0];
  assign mem_202_5_W0_clk = W0_clk;
  assign mem_202_5_W0_data = W0_data[47:40];
  assign mem_202_5_W0_en = W0_en & W0_addr_sel == 8'hca;
  assign mem_202_5_W0_mask = W0_mask[5];
  assign mem_202_6_R0_addr = R0_addr[25:0];
  assign mem_202_6_R0_clk = R0_clk;
  assign mem_202_6_R0_en = R0_en & R0_addr_sel == 8'hca;
  assign mem_202_6_W0_addr = W0_addr[25:0];
  assign mem_202_6_W0_clk = W0_clk;
  assign mem_202_6_W0_data = W0_data[55:48];
  assign mem_202_6_W0_en = W0_en & W0_addr_sel == 8'hca;
  assign mem_202_6_W0_mask = W0_mask[6];
  assign mem_202_7_R0_addr = R0_addr[25:0];
  assign mem_202_7_R0_clk = R0_clk;
  assign mem_202_7_R0_en = R0_en & R0_addr_sel == 8'hca;
  assign mem_202_7_W0_addr = W0_addr[25:0];
  assign mem_202_7_W0_clk = W0_clk;
  assign mem_202_7_W0_data = W0_data[63:56];
  assign mem_202_7_W0_en = W0_en & W0_addr_sel == 8'hca;
  assign mem_202_7_W0_mask = W0_mask[7];
  assign mem_203_0_R0_addr = R0_addr[25:0];
  assign mem_203_0_R0_clk = R0_clk;
  assign mem_203_0_R0_en = R0_en & R0_addr_sel == 8'hcb;
  assign mem_203_0_W0_addr = W0_addr[25:0];
  assign mem_203_0_W0_clk = W0_clk;
  assign mem_203_0_W0_data = W0_data[7:0];
  assign mem_203_0_W0_en = W0_en & W0_addr_sel == 8'hcb;
  assign mem_203_0_W0_mask = W0_mask[0];
  assign mem_203_1_R0_addr = R0_addr[25:0];
  assign mem_203_1_R0_clk = R0_clk;
  assign mem_203_1_R0_en = R0_en & R0_addr_sel == 8'hcb;
  assign mem_203_1_W0_addr = W0_addr[25:0];
  assign mem_203_1_W0_clk = W0_clk;
  assign mem_203_1_W0_data = W0_data[15:8];
  assign mem_203_1_W0_en = W0_en & W0_addr_sel == 8'hcb;
  assign mem_203_1_W0_mask = W0_mask[1];
  assign mem_203_2_R0_addr = R0_addr[25:0];
  assign mem_203_2_R0_clk = R0_clk;
  assign mem_203_2_R0_en = R0_en & R0_addr_sel == 8'hcb;
  assign mem_203_2_W0_addr = W0_addr[25:0];
  assign mem_203_2_W0_clk = W0_clk;
  assign mem_203_2_W0_data = W0_data[23:16];
  assign mem_203_2_W0_en = W0_en & W0_addr_sel == 8'hcb;
  assign mem_203_2_W0_mask = W0_mask[2];
  assign mem_203_3_R0_addr = R0_addr[25:0];
  assign mem_203_3_R0_clk = R0_clk;
  assign mem_203_3_R0_en = R0_en & R0_addr_sel == 8'hcb;
  assign mem_203_3_W0_addr = W0_addr[25:0];
  assign mem_203_3_W0_clk = W0_clk;
  assign mem_203_3_W0_data = W0_data[31:24];
  assign mem_203_3_W0_en = W0_en & W0_addr_sel == 8'hcb;
  assign mem_203_3_W0_mask = W0_mask[3];
  assign mem_203_4_R0_addr = R0_addr[25:0];
  assign mem_203_4_R0_clk = R0_clk;
  assign mem_203_4_R0_en = R0_en & R0_addr_sel == 8'hcb;
  assign mem_203_4_W0_addr = W0_addr[25:0];
  assign mem_203_4_W0_clk = W0_clk;
  assign mem_203_4_W0_data = W0_data[39:32];
  assign mem_203_4_W0_en = W0_en & W0_addr_sel == 8'hcb;
  assign mem_203_4_W0_mask = W0_mask[4];
  assign mem_203_5_R0_addr = R0_addr[25:0];
  assign mem_203_5_R0_clk = R0_clk;
  assign mem_203_5_R0_en = R0_en & R0_addr_sel == 8'hcb;
  assign mem_203_5_W0_addr = W0_addr[25:0];
  assign mem_203_5_W0_clk = W0_clk;
  assign mem_203_5_W0_data = W0_data[47:40];
  assign mem_203_5_W0_en = W0_en & W0_addr_sel == 8'hcb;
  assign mem_203_5_W0_mask = W0_mask[5];
  assign mem_203_6_R0_addr = R0_addr[25:0];
  assign mem_203_6_R0_clk = R0_clk;
  assign mem_203_6_R0_en = R0_en & R0_addr_sel == 8'hcb;
  assign mem_203_6_W0_addr = W0_addr[25:0];
  assign mem_203_6_W0_clk = W0_clk;
  assign mem_203_6_W0_data = W0_data[55:48];
  assign mem_203_6_W0_en = W0_en & W0_addr_sel == 8'hcb;
  assign mem_203_6_W0_mask = W0_mask[6];
  assign mem_203_7_R0_addr = R0_addr[25:0];
  assign mem_203_7_R0_clk = R0_clk;
  assign mem_203_7_R0_en = R0_en & R0_addr_sel == 8'hcb;
  assign mem_203_7_W0_addr = W0_addr[25:0];
  assign mem_203_7_W0_clk = W0_clk;
  assign mem_203_7_W0_data = W0_data[63:56];
  assign mem_203_7_W0_en = W0_en & W0_addr_sel == 8'hcb;
  assign mem_203_7_W0_mask = W0_mask[7];
  assign mem_204_0_R0_addr = R0_addr[25:0];
  assign mem_204_0_R0_clk = R0_clk;
  assign mem_204_0_R0_en = R0_en & R0_addr_sel == 8'hcc;
  assign mem_204_0_W0_addr = W0_addr[25:0];
  assign mem_204_0_W0_clk = W0_clk;
  assign mem_204_0_W0_data = W0_data[7:0];
  assign mem_204_0_W0_en = W0_en & W0_addr_sel == 8'hcc;
  assign mem_204_0_W0_mask = W0_mask[0];
  assign mem_204_1_R0_addr = R0_addr[25:0];
  assign mem_204_1_R0_clk = R0_clk;
  assign mem_204_1_R0_en = R0_en & R0_addr_sel == 8'hcc;
  assign mem_204_1_W0_addr = W0_addr[25:0];
  assign mem_204_1_W0_clk = W0_clk;
  assign mem_204_1_W0_data = W0_data[15:8];
  assign mem_204_1_W0_en = W0_en & W0_addr_sel == 8'hcc;
  assign mem_204_1_W0_mask = W0_mask[1];
  assign mem_204_2_R0_addr = R0_addr[25:0];
  assign mem_204_2_R0_clk = R0_clk;
  assign mem_204_2_R0_en = R0_en & R0_addr_sel == 8'hcc;
  assign mem_204_2_W0_addr = W0_addr[25:0];
  assign mem_204_2_W0_clk = W0_clk;
  assign mem_204_2_W0_data = W0_data[23:16];
  assign mem_204_2_W0_en = W0_en & W0_addr_sel == 8'hcc;
  assign mem_204_2_W0_mask = W0_mask[2];
  assign mem_204_3_R0_addr = R0_addr[25:0];
  assign mem_204_3_R0_clk = R0_clk;
  assign mem_204_3_R0_en = R0_en & R0_addr_sel == 8'hcc;
  assign mem_204_3_W0_addr = W0_addr[25:0];
  assign mem_204_3_W0_clk = W0_clk;
  assign mem_204_3_W0_data = W0_data[31:24];
  assign mem_204_3_W0_en = W0_en & W0_addr_sel == 8'hcc;
  assign mem_204_3_W0_mask = W0_mask[3];
  assign mem_204_4_R0_addr = R0_addr[25:0];
  assign mem_204_4_R0_clk = R0_clk;
  assign mem_204_4_R0_en = R0_en & R0_addr_sel == 8'hcc;
  assign mem_204_4_W0_addr = W0_addr[25:0];
  assign mem_204_4_W0_clk = W0_clk;
  assign mem_204_4_W0_data = W0_data[39:32];
  assign mem_204_4_W0_en = W0_en & W0_addr_sel == 8'hcc;
  assign mem_204_4_W0_mask = W0_mask[4];
  assign mem_204_5_R0_addr = R0_addr[25:0];
  assign mem_204_5_R0_clk = R0_clk;
  assign mem_204_5_R0_en = R0_en & R0_addr_sel == 8'hcc;
  assign mem_204_5_W0_addr = W0_addr[25:0];
  assign mem_204_5_W0_clk = W0_clk;
  assign mem_204_5_W0_data = W0_data[47:40];
  assign mem_204_5_W0_en = W0_en & W0_addr_sel == 8'hcc;
  assign mem_204_5_W0_mask = W0_mask[5];
  assign mem_204_6_R0_addr = R0_addr[25:0];
  assign mem_204_6_R0_clk = R0_clk;
  assign mem_204_6_R0_en = R0_en & R0_addr_sel == 8'hcc;
  assign mem_204_6_W0_addr = W0_addr[25:0];
  assign mem_204_6_W0_clk = W0_clk;
  assign mem_204_6_W0_data = W0_data[55:48];
  assign mem_204_6_W0_en = W0_en & W0_addr_sel == 8'hcc;
  assign mem_204_6_W0_mask = W0_mask[6];
  assign mem_204_7_R0_addr = R0_addr[25:0];
  assign mem_204_7_R0_clk = R0_clk;
  assign mem_204_7_R0_en = R0_en & R0_addr_sel == 8'hcc;
  assign mem_204_7_W0_addr = W0_addr[25:0];
  assign mem_204_7_W0_clk = W0_clk;
  assign mem_204_7_W0_data = W0_data[63:56];
  assign mem_204_7_W0_en = W0_en & W0_addr_sel == 8'hcc;
  assign mem_204_7_W0_mask = W0_mask[7];
  assign mem_205_0_R0_addr = R0_addr[25:0];
  assign mem_205_0_R0_clk = R0_clk;
  assign mem_205_0_R0_en = R0_en & R0_addr_sel == 8'hcd;
  assign mem_205_0_W0_addr = W0_addr[25:0];
  assign mem_205_0_W0_clk = W0_clk;
  assign mem_205_0_W0_data = W0_data[7:0];
  assign mem_205_0_W0_en = W0_en & W0_addr_sel == 8'hcd;
  assign mem_205_0_W0_mask = W0_mask[0];
  assign mem_205_1_R0_addr = R0_addr[25:0];
  assign mem_205_1_R0_clk = R0_clk;
  assign mem_205_1_R0_en = R0_en & R0_addr_sel == 8'hcd;
  assign mem_205_1_W0_addr = W0_addr[25:0];
  assign mem_205_1_W0_clk = W0_clk;
  assign mem_205_1_W0_data = W0_data[15:8];
  assign mem_205_1_W0_en = W0_en & W0_addr_sel == 8'hcd;
  assign mem_205_1_W0_mask = W0_mask[1];
  assign mem_205_2_R0_addr = R0_addr[25:0];
  assign mem_205_2_R0_clk = R0_clk;
  assign mem_205_2_R0_en = R0_en & R0_addr_sel == 8'hcd;
  assign mem_205_2_W0_addr = W0_addr[25:0];
  assign mem_205_2_W0_clk = W0_clk;
  assign mem_205_2_W0_data = W0_data[23:16];
  assign mem_205_2_W0_en = W0_en & W0_addr_sel == 8'hcd;
  assign mem_205_2_W0_mask = W0_mask[2];
  assign mem_205_3_R0_addr = R0_addr[25:0];
  assign mem_205_3_R0_clk = R0_clk;
  assign mem_205_3_R0_en = R0_en & R0_addr_sel == 8'hcd;
  assign mem_205_3_W0_addr = W0_addr[25:0];
  assign mem_205_3_W0_clk = W0_clk;
  assign mem_205_3_W0_data = W0_data[31:24];
  assign mem_205_3_W0_en = W0_en & W0_addr_sel == 8'hcd;
  assign mem_205_3_W0_mask = W0_mask[3];
  assign mem_205_4_R0_addr = R0_addr[25:0];
  assign mem_205_4_R0_clk = R0_clk;
  assign mem_205_4_R0_en = R0_en & R0_addr_sel == 8'hcd;
  assign mem_205_4_W0_addr = W0_addr[25:0];
  assign mem_205_4_W0_clk = W0_clk;
  assign mem_205_4_W0_data = W0_data[39:32];
  assign mem_205_4_W0_en = W0_en & W0_addr_sel == 8'hcd;
  assign mem_205_4_W0_mask = W0_mask[4];
  assign mem_205_5_R0_addr = R0_addr[25:0];
  assign mem_205_5_R0_clk = R0_clk;
  assign mem_205_5_R0_en = R0_en & R0_addr_sel == 8'hcd;
  assign mem_205_5_W0_addr = W0_addr[25:0];
  assign mem_205_5_W0_clk = W0_clk;
  assign mem_205_5_W0_data = W0_data[47:40];
  assign mem_205_5_W0_en = W0_en & W0_addr_sel == 8'hcd;
  assign mem_205_5_W0_mask = W0_mask[5];
  assign mem_205_6_R0_addr = R0_addr[25:0];
  assign mem_205_6_R0_clk = R0_clk;
  assign mem_205_6_R0_en = R0_en & R0_addr_sel == 8'hcd;
  assign mem_205_6_W0_addr = W0_addr[25:0];
  assign mem_205_6_W0_clk = W0_clk;
  assign mem_205_6_W0_data = W0_data[55:48];
  assign mem_205_6_W0_en = W0_en & W0_addr_sel == 8'hcd;
  assign mem_205_6_W0_mask = W0_mask[6];
  assign mem_205_7_R0_addr = R0_addr[25:0];
  assign mem_205_7_R0_clk = R0_clk;
  assign mem_205_7_R0_en = R0_en & R0_addr_sel == 8'hcd;
  assign mem_205_7_W0_addr = W0_addr[25:0];
  assign mem_205_7_W0_clk = W0_clk;
  assign mem_205_7_W0_data = W0_data[63:56];
  assign mem_205_7_W0_en = W0_en & W0_addr_sel == 8'hcd;
  assign mem_205_7_W0_mask = W0_mask[7];
  assign mem_206_0_R0_addr = R0_addr[25:0];
  assign mem_206_0_R0_clk = R0_clk;
  assign mem_206_0_R0_en = R0_en & R0_addr_sel == 8'hce;
  assign mem_206_0_W0_addr = W0_addr[25:0];
  assign mem_206_0_W0_clk = W0_clk;
  assign mem_206_0_W0_data = W0_data[7:0];
  assign mem_206_0_W0_en = W0_en & W0_addr_sel == 8'hce;
  assign mem_206_0_W0_mask = W0_mask[0];
  assign mem_206_1_R0_addr = R0_addr[25:0];
  assign mem_206_1_R0_clk = R0_clk;
  assign mem_206_1_R0_en = R0_en & R0_addr_sel == 8'hce;
  assign mem_206_1_W0_addr = W0_addr[25:0];
  assign mem_206_1_W0_clk = W0_clk;
  assign mem_206_1_W0_data = W0_data[15:8];
  assign mem_206_1_W0_en = W0_en & W0_addr_sel == 8'hce;
  assign mem_206_1_W0_mask = W0_mask[1];
  assign mem_206_2_R0_addr = R0_addr[25:0];
  assign mem_206_2_R0_clk = R0_clk;
  assign mem_206_2_R0_en = R0_en & R0_addr_sel == 8'hce;
  assign mem_206_2_W0_addr = W0_addr[25:0];
  assign mem_206_2_W0_clk = W0_clk;
  assign mem_206_2_W0_data = W0_data[23:16];
  assign mem_206_2_W0_en = W0_en & W0_addr_sel == 8'hce;
  assign mem_206_2_W0_mask = W0_mask[2];
  assign mem_206_3_R0_addr = R0_addr[25:0];
  assign mem_206_3_R0_clk = R0_clk;
  assign mem_206_3_R0_en = R0_en & R0_addr_sel == 8'hce;
  assign mem_206_3_W0_addr = W0_addr[25:0];
  assign mem_206_3_W0_clk = W0_clk;
  assign mem_206_3_W0_data = W0_data[31:24];
  assign mem_206_3_W0_en = W0_en & W0_addr_sel == 8'hce;
  assign mem_206_3_W0_mask = W0_mask[3];
  assign mem_206_4_R0_addr = R0_addr[25:0];
  assign mem_206_4_R0_clk = R0_clk;
  assign mem_206_4_R0_en = R0_en & R0_addr_sel == 8'hce;
  assign mem_206_4_W0_addr = W0_addr[25:0];
  assign mem_206_4_W0_clk = W0_clk;
  assign mem_206_4_W0_data = W0_data[39:32];
  assign mem_206_4_W0_en = W0_en & W0_addr_sel == 8'hce;
  assign mem_206_4_W0_mask = W0_mask[4];
  assign mem_206_5_R0_addr = R0_addr[25:0];
  assign mem_206_5_R0_clk = R0_clk;
  assign mem_206_5_R0_en = R0_en & R0_addr_sel == 8'hce;
  assign mem_206_5_W0_addr = W0_addr[25:0];
  assign mem_206_5_W0_clk = W0_clk;
  assign mem_206_5_W0_data = W0_data[47:40];
  assign mem_206_5_W0_en = W0_en & W0_addr_sel == 8'hce;
  assign mem_206_5_W0_mask = W0_mask[5];
  assign mem_206_6_R0_addr = R0_addr[25:0];
  assign mem_206_6_R0_clk = R0_clk;
  assign mem_206_6_R0_en = R0_en & R0_addr_sel == 8'hce;
  assign mem_206_6_W0_addr = W0_addr[25:0];
  assign mem_206_6_W0_clk = W0_clk;
  assign mem_206_6_W0_data = W0_data[55:48];
  assign mem_206_6_W0_en = W0_en & W0_addr_sel == 8'hce;
  assign mem_206_6_W0_mask = W0_mask[6];
  assign mem_206_7_R0_addr = R0_addr[25:0];
  assign mem_206_7_R0_clk = R0_clk;
  assign mem_206_7_R0_en = R0_en & R0_addr_sel == 8'hce;
  assign mem_206_7_W0_addr = W0_addr[25:0];
  assign mem_206_7_W0_clk = W0_clk;
  assign mem_206_7_W0_data = W0_data[63:56];
  assign mem_206_7_W0_en = W0_en & W0_addr_sel == 8'hce;
  assign mem_206_7_W0_mask = W0_mask[7];
  assign mem_207_0_R0_addr = R0_addr[25:0];
  assign mem_207_0_R0_clk = R0_clk;
  assign mem_207_0_R0_en = R0_en & R0_addr_sel == 8'hcf;
  assign mem_207_0_W0_addr = W0_addr[25:0];
  assign mem_207_0_W0_clk = W0_clk;
  assign mem_207_0_W0_data = W0_data[7:0];
  assign mem_207_0_W0_en = W0_en & W0_addr_sel == 8'hcf;
  assign mem_207_0_W0_mask = W0_mask[0];
  assign mem_207_1_R0_addr = R0_addr[25:0];
  assign mem_207_1_R0_clk = R0_clk;
  assign mem_207_1_R0_en = R0_en & R0_addr_sel == 8'hcf;
  assign mem_207_1_W0_addr = W0_addr[25:0];
  assign mem_207_1_W0_clk = W0_clk;
  assign mem_207_1_W0_data = W0_data[15:8];
  assign mem_207_1_W0_en = W0_en & W0_addr_sel == 8'hcf;
  assign mem_207_1_W0_mask = W0_mask[1];
  assign mem_207_2_R0_addr = R0_addr[25:0];
  assign mem_207_2_R0_clk = R0_clk;
  assign mem_207_2_R0_en = R0_en & R0_addr_sel == 8'hcf;
  assign mem_207_2_W0_addr = W0_addr[25:0];
  assign mem_207_2_W0_clk = W0_clk;
  assign mem_207_2_W0_data = W0_data[23:16];
  assign mem_207_2_W0_en = W0_en & W0_addr_sel == 8'hcf;
  assign mem_207_2_W0_mask = W0_mask[2];
  assign mem_207_3_R0_addr = R0_addr[25:0];
  assign mem_207_3_R0_clk = R0_clk;
  assign mem_207_3_R0_en = R0_en & R0_addr_sel == 8'hcf;
  assign mem_207_3_W0_addr = W0_addr[25:0];
  assign mem_207_3_W0_clk = W0_clk;
  assign mem_207_3_W0_data = W0_data[31:24];
  assign mem_207_3_W0_en = W0_en & W0_addr_sel == 8'hcf;
  assign mem_207_3_W0_mask = W0_mask[3];
  assign mem_207_4_R0_addr = R0_addr[25:0];
  assign mem_207_4_R0_clk = R0_clk;
  assign mem_207_4_R0_en = R0_en & R0_addr_sel == 8'hcf;
  assign mem_207_4_W0_addr = W0_addr[25:0];
  assign mem_207_4_W0_clk = W0_clk;
  assign mem_207_4_W0_data = W0_data[39:32];
  assign mem_207_4_W0_en = W0_en & W0_addr_sel == 8'hcf;
  assign mem_207_4_W0_mask = W0_mask[4];
  assign mem_207_5_R0_addr = R0_addr[25:0];
  assign mem_207_5_R0_clk = R0_clk;
  assign mem_207_5_R0_en = R0_en & R0_addr_sel == 8'hcf;
  assign mem_207_5_W0_addr = W0_addr[25:0];
  assign mem_207_5_W0_clk = W0_clk;
  assign mem_207_5_W0_data = W0_data[47:40];
  assign mem_207_5_W0_en = W0_en & W0_addr_sel == 8'hcf;
  assign mem_207_5_W0_mask = W0_mask[5];
  assign mem_207_6_R0_addr = R0_addr[25:0];
  assign mem_207_6_R0_clk = R0_clk;
  assign mem_207_6_R0_en = R0_en & R0_addr_sel == 8'hcf;
  assign mem_207_6_W0_addr = W0_addr[25:0];
  assign mem_207_6_W0_clk = W0_clk;
  assign mem_207_6_W0_data = W0_data[55:48];
  assign mem_207_6_W0_en = W0_en & W0_addr_sel == 8'hcf;
  assign mem_207_6_W0_mask = W0_mask[6];
  assign mem_207_7_R0_addr = R0_addr[25:0];
  assign mem_207_7_R0_clk = R0_clk;
  assign mem_207_7_R0_en = R0_en & R0_addr_sel == 8'hcf;
  assign mem_207_7_W0_addr = W0_addr[25:0];
  assign mem_207_7_W0_clk = W0_clk;
  assign mem_207_7_W0_data = W0_data[63:56];
  assign mem_207_7_W0_en = W0_en & W0_addr_sel == 8'hcf;
  assign mem_207_7_W0_mask = W0_mask[7];
  assign mem_208_0_R0_addr = R0_addr[25:0];
  assign mem_208_0_R0_clk = R0_clk;
  assign mem_208_0_R0_en = R0_en & R0_addr_sel == 8'hd0;
  assign mem_208_0_W0_addr = W0_addr[25:0];
  assign mem_208_0_W0_clk = W0_clk;
  assign mem_208_0_W0_data = W0_data[7:0];
  assign mem_208_0_W0_en = W0_en & W0_addr_sel == 8'hd0;
  assign mem_208_0_W0_mask = W0_mask[0];
  assign mem_208_1_R0_addr = R0_addr[25:0];
  assign mem_208_1_R0_clk = R0_clk;
  assign mem_208_1_R0_en = R0_en & R0_addr_sel == 8'hd0;
  assign mem_208_1_W0_addr = W0_addr[25:0];
  assign mem_208_1_W0_clk = W0_clk;
  assign mem_208_1_W0_data = W0_data[15:8];
  assign mem_208_1_W0_en = W0_en & W0_addr_sel == 8'hd0;
  assign mem_208_1_W0_mask = W0_mask[1];
  assign mem_208_2_R0_addr = R0_addr[25:0];
  assign mem_208_2_R0_clk = R0_clk;
  assign mem_208_2_R0_en = R0_en & R0_addr_sel == 8'hd0;
  assign mem_208_2_W0_addr = W0_addr[25:0];
  assign mem_208_2_W0_clk = W0_clk;
  assign mem_208_2_W0_data = W0_data[23:16];
  assign mem_208_2_W0_en = W0_en & W0_addr_sel == 8'hd0;
  assign mem_208_2_W0_mask = W0_mask[2];
  assign mem_208_3_R0_addr = R0_addr[25:0];
  assign mem_208_3_R0_clk = R0_clk;
  assign mem_208_3_R0_en = R0_en & R0_addr_sel == 8'hd0;
  assign mem_208_3_W0_addr = W0_addr[25:0];
  assign mem_208_3_W0_clk = W0_clk;
  assign mem_208_3_W0_data = W0_data[31:24];
  assign mem_208_3_W0_en = W0_en & W0_addr_sel == 8'hd0;
  assign mem_208_3_W0_mask = W0_mask[3];
  assign mem_208_4_R0_addr = R0_addr[25:0];
  assign mem_208_4_R0_clk = R0_clk;
  assign mem_208_4_R0_en = R0_en & R0_addr_sel == 8'hd0;
  assign mem_208_4_W0_addr = W0_addr[25:0];
  assign mem_208_4_W0_clk = W0_clk;
  assign mem_208_4_W0_data = W0_data[39:32];
  assign mem_208_4_W0_en = W0_en & W0_addr_sel == 8'hd0;
  assign mem_208_4_W0_mask = W0_mask[4];
  assign mem_208_5_R0_addr = R0_addr[25:0];
  assign mem_208_5_R0_clk = R0_clk;
  assign mem_208_5_R0_en = R0_en & R0_addr_sel == 8'hd0;
  assign mem_208_5_W0_addr = W0_addr[25:0];
  assign mem_208_5_W0_clk = W0_clk;
  assign mem_208_5_W0_data = W0_data[47:40];
  assign mem_208_5_W0_en = W0_en & W0_addr_sel == 8'hd0;
  assign mem_208_5_W0_mask = W0_mask[5];
  assign mem_208_6_R0_addr = R0_addr[25:0];
  assign mem_208_6_R0_clk = R0_clk;
  assign mem_208_6_R0_en = R0_en & R0_addr_sel == 8'hd0;
  assign mem_208_6_W0_addr = W0_addr[25:0];
  assign mem_208_6_W0_clk = W0_clk;
  assign mem_208_6_W0_data = W0_data[55:48];
  assign mem_208_6_W0_en = W0_en & W0_addr_sel == 8'hd0;
  assign mem_208_6_W0_mask = W0_mask[6];
  assign mem_208_7_R0_addr = R0_addr[25:0];
  assign mem_208_7_R0_clk = R0_clk;
  assign mem_208_7_R0_en = R0_en & R0_addr_sel == 8'hd0;
  assign mem_208_7_W0_addr = W0_addr[25:0];
  assign mem_208_7_W0_clk = W0_clk;
  assign mem_208_7_W0_data = W0_data[63:56];
  assign mem_208_7_W0_en = W0_en & W0_addr_sel == 8'hd0;
  assign mem_208_7_W0_mask = W0_mask[7];
  assign mem_209_0_R0_addr = R0_addr[25:0];
  assign mem_209_0_R0_clk = R0_clk;
  assign mem_209_0_R0_en = R0_en & R0_addr_sel == 8'hd1;
  assign mem_209_0_W0_addr = W0_addr[25:0];
  assign mem_209_0_W0_clk = W0_clk;
  assign mem_209_0_W0_data = W0_data[7:0];
  assign mem_209_0_W0_en = W0_en & W0_addr_sel == 8'hd1;
  assign mem_209_0_W0_mask = W0_mask[0];
  assign mem_209_1_R0_addr = R0_addr[25:0];
  assign mem_209_1_R0_clk = R0_clk;
  assign mem_209_1_R0_en = R0_en & R0_addr_sel == 8'hd1;
  assign mem_209_1_W0_addr = W0_addr[25:0];
  assign mem_209_1_W0_clk = W0_clk;
  assign mem_209_1_W0_data = W0_data[15:8];
  assign mem_209_1_W0_en = W0_en & W0_addr_sel == 8'hd1;
  assign mem_209_1_W0_mask = W0_mask[1];
  assign mem_209_2_R0_addr = R0_addr[25:0];
  assign mem_209_2_R0_clk = R0_clk;
  assign mem_209_2_R0_en = R0_en & R0_addr_sel == 8'hd1;
  assign mem_209_2_W0_addr = W0_addr[25:0];
  assign mem_209_2_W0_clk = W0_clk;
  assign mem_209_2_W0_data = W0_data[23:16];
  assign mem_209_2_W0_en = W0_en & W0_addr_sel == 8'hd1;
  assign mem_209_2_W0_mask = W0_mask[2];
  assign mem_209_3_R0_addr = R0_addr[25:0];
  assign mem_209_3_R0_clk = R0_clk;
  assign mem_209_3_R0_en = R0_en & R0_addr_sel == 8'hd1;
  assign mem_209_3_W0_addr = W0_addr[25:0];
  assign mem_209_3_W0_clk = W0_clk;
  assign mem_209_3_W0_data = W0_data[31:24];
  assign mem_209_3_W0_en = W0_en & W0_addr_sel == 8'hd1;
  assign mem_209_3_W0_mask = W0_mask[3];
  assign mem_209_4_R0_addr = R0_addr[25:0];
  assign mem_209_4_R0_clk = R0_clk;
  assign mem_209_4_R0_en = R0_en & R0_addr_sel == 8'hd1;
  assign mem_209_4_W0_addr = W0_addr[25:0];
  assign mem_209_4_W0_clk = W0_clk;
  assign mem_209_4_W0_data = W0_data[39:32];
  assign mem_209_4_W0_en = W0_en & W0_addr_sel == 8'hd1;
  assign mem_209_4_W0_mask = W0_mask[4];
  assign mem_209_5_R0_addr = R0_addr[25:0];
  assign mem_209_5_R0_clk = R0_clk;
  assign mem_209_5_R0_en = R0_en & R0_addr_sel == 8'hd1;
  assign mem_209_5_W0_addr = W0_addr[25:0];
  assign mem_209_5_W0_clk = W0_clk;
  assign mem_209_5_W0_data = W0_data[47:40];
  assign mem_209_5_W0_en = W0_en & W0_addr_sel == 8'hd1;
  assign mem_209_5_W0_mask = W0_mask[5];
  assign mem_209_6_R0_addr = R0_addr[25:0];
  assign mem_209_6_R0_clk = R0_clk;
  assign mem_209_6_R0_en = R0_en & R0_addr_sel == 8'hd1;
  assign mem_209_6_W0_addr = W0_addr[25:0];
  assign mem_209_6_W0_clk = W0_clk;
  assign mem_209_6_W0_data = W0_data[55:48];
  assign mem_209_6_W0_en = W0_en & W0_addr_sel == 8'hd1;
  assign mem_209_6_W0_mask = W0_mask[6];
  assign mem_209_7_R0_addr = R0_addr[25:0];
  assign mem_209_7_R0_clk = R0_clk;
  assign mem_209_7_R0_en = R0_en & R0_addr_sel == 8'hd1;
  assign mem_209_7_W0_addr = W0_addr[25:0];
  assign mem_209_7_W0_clk = W0_clk;
  assign mem_209_7_W0_data = W0_data[63:56];
  assign mem_209_7_W0_en = W0_en & W0_addr_sel == 8'hd1;
  assign mem_209_7_W0_mask = W0_mask[7];
  assign mem_210_0_R0_addr = R0_addr[25:0];
  assign mem_210_0_R0_clk = R0_clk;
  assign mem_210_0_R0_en = R0_en & R0_addr_sel == 8'hd2;
  assign mem_210_0_W0_addr = W0_addr[25:0];
  assign mem_210_0_W0_clk = W0_clk;
  assign mem_210_0_W0_data = W0_data[7:0];
  assign mem_210_0_W0_en = W0_en & W0_addr_sel == 8'hd2;
  assign mem_210_0_W0_mask = W0_mask[0];
  assign mem_210_1_R0_addr = R0_addr[25:0];
  assign mem_210_1_R0_clk = R0_clk;
  assign mem_210_1_R0_en = R0_en & R0_addr_sel == 8'hd2;
  assign mem_210_1_W0_addr = W0_addr[25:0];
  assign mem_210_1_W0_clk = W0_clk;
  assign mem_210_1_W0_data = W0_data[15:8];
  assign mem_210_1_W0_en = W0_en & W0_addr_sel == 8'hd2;
  assign mem_210_1_W0_mask = W0_mask[1];
  assign mem_210_2_R0_addr = R0_addr[25:0];
  assign mem_210_2_R0_clk = R0_clk;
  assign mem_210_2_R0_en = R0_en & R0_addr_sel == 8'hd2;
  assign mem_210_2_W0_addr = W0_addr[25:0];
  assign mem_210_2_W0_clk = W0_clk;
  assign mem_210_2_W0_data = W0_data[23:16];
  assign mem_210_2_W0_en = W0_en & W0_addr_sel == 8'hd2;
  assign mem_210_2_W0_mask = W0_mask[2];
  assign mem_210_3_R0_addr = R0_addr[25:0];
  assign mem_210_3_R0_clk = R0_clk;
  assign mem_210_3_R0_en = R0_en & R0_addr_sel == 8'hd2;
  assign mem_210_3_W0_addr = W0_addr[25:0];
  assign mem_210_3_W0_clk = W0_clk;
  assign mem_210_3_W0_data = W0_data[31:24];
  assign mem_210_3_W0_en = W0_en & W0_addr_sel == 8'hd2;
  assign mem_210_3_W0_mask = W0_mask[3];
  assign mem_210_4_R0_addr = R0_addr[25:0];
  assign mem_210_4_R0_clk = R0_clk;
  assign mem_210_4_R0_en = R0_en & R0_addr_sel == 8'hd2;
  assign mem_210_4_W0_addr = W0_addr[25:0];
  assign mem_210_4_W0_clk = W0_clk;
  assign mem_210_4_W0_data = W0_data[39:32];
  assign mem_210_4_W0_en = W0_en & W0_addr_sel == 8'hd2;
  assign mem_210_4_W0_mask = W0_mask[4];
  assign mem_210_5_R0_addr = R0_addr[25:0];
  assign mem_210_5_R0_clk = R0_clk;
  assign mem_210_5_R0_en = R0_en & R0_addr_sel == 8'hd2;
  assign mem_210_5_W0_addr = W0_addr[25:0];
  assign mem_210_5_W0_clk = W0_clk;
  assign mem_210_5_W0_data = W0_data[47:40];
  assign mem_210_5_W0_en = W0_en & W0_addr_sel == 8'hd2;
  assign mem_210_5_W0_mask = W0_mask[5];
  assign mem_210_6_R0_addr = R0_addr[25:0];
  assign mem_210_6_R0_clk = R0_clk;
  assign mem_210_6_R0_en = R0_en & R0_addr_sel == 8'hd2;
  assign mem_210_6_W0_addr = W0_addr[25:0];
  assign mem_210_6_W0_clk = W0_clk;
  assign mem_210_6_W0_data = W0_data[55:48];
  assign mem_210_6_W0_en = W0_en & W0_addr_sel == 8'hd2;
  assign mem_210_6_W0_mask = W0_mask[6];
  assign mem_210_7_R0_addr = R0_addr[25:0];
  assign mem_210_7_R0_clk = R0_clk;
  assign mem_210_7_R0_en = R0_en & R0_addr_sel == 8'hd2;
  assign mem_210_7_W0_addr = W0_addr[25:0];
  assign mem_210_7_W0_clk = W0_clk;
  assign mem_210_7_W0_data = W0_data[63:56];
  assign mem_210_7_W0_en = W0_en & W0_addr_sel == 8'hd2;
  assign mem_210_7_W0_mask = W0_mask[7];
  assign mem_211_0_R0_addr = R0_addr[25:0];
  assign mem_211_0_R0_clk = R0_clk;
  assign mem_211_0_R0_en = R0_en & R0_addr_sel == 8'hd3;
  assign mem_211_0_W0_addr = W0_addr[25:0];
  assign mem_211_0_W0_clk = W0_clk;
  assign mem_211_0_W0_data = W0_data[7:0];
  assign mem_211_0_W0_en = W0_en & W0_addr_sel == 8'hd3;
  assign mem_211_0_W0_mask = W0_mask[0];
  assign mem_211_1_R0_addr = R0_addr[25:0];
  assign mem_211_1_R0_clk = R0_clk;
  assign mem_211_1_R0_en = R0_en & R0_addr_sel == 8'hd3;
  assign mem_211_1_W0_addr = W0_addr[25:0];
  assign mem_211_1_W0_clk = W0_clk;
  assign mem_211_1_W0_data = W0_data[15:8];
  assign mem_211_1_W0_en = W0_en & W0_addr_sel == 8'hd3;
  assign mem_211_1_W0_mask = W0_mask[1];
  assign mem_211_2_R0_addr = R0_addr[25:0];
  assign mem_211_2_R0_clk = R0_clk;
  assign mem_211_2_R0_en = R0_en & R0_addr_sel == 8'hd3;
  assign mem_211_2_W0_addr = W0_addr[25:0];
  assign mem_211_2_W0_clk = W0_clk;
  assign mem_211_2_W0_data = W0_data[23:16];
  assign mem_211_2_W0_en = W0_en & W0_addr_sel == 8'hd3;
  assign mem_211_2_W0_mask = W0_mask[2];
  assign mem_211_3_R0_addr = R0_addr[25:0];
  assign mem_211_3_R0_clk = R0_clk;
  assign mem_211_3_R0_en = R0_en & R0_addr_sel == 8'hd3;
  assign mem_211_3_W0_addr = W0_addr[25:0];
  assign mem_211_3_W0_clk = W0_clk;
  assign mem_211_3_W0_data = W0_data[31:24];
  assign mem_211_3_W0_en = W0_en & W0_addr_sel == 8'hd3;
  assign mem_211_3_W0_mask = W0_mask[3];
  assign mem_211_4_R0_addr = R0_addr[25:0];
  assign mem_211_4_R0_clk = R0_clk;
  assign mem_211_4_R0_en = R0_en & R0_addr_sel == 8'hd3;
  assign mem_211_4_W0_addr = W0_addr[25:0];
  assign mem_211_4_W0_clk = W0_clk;
  assign mem_211_4_W0_data = W0_data[39:32];
  assign mem_211_4_W0_en = W0_en & W0_addr_sel == 8'hd3;
  assign mem_211_4_W0_mask = W0_mask[4];
  assign mem_211_5_R0_addr = R0_addr[25:0];
  assign mem_211_5_R0_clk = R0_clk;
  assign mem_211_5_R0_en = R0_en & R0_addr_sel == 8'hd3;
  assign mem_211_5_W0_addr = W0_addr[25:0];
  assign mem_211_5_W0_clk = W0_clk;
  assign mem_211_5_W0_data = W0_data[47:40];
  assign mem_211_5_W0_en = W0_en & W0_addr_sel == 8'hd3;
  assign mem_211_5_W0_mask = W0_mask[5];
  assign mem_211_6_R0_addr = R0_addr[25:0];
  assign mem_211_6_R0_clk = R0_clk;
  assign mem_211_6_R0_en = R0_en & R0_addr_sel == 8'hd3;
  assign mem_211_6_W0_addr = W0_addr[25:0];
  assign mem_211_6_W0_clk = W0_clk;
  assign mem_211_6_W0_data = W0_data[55:48];
  assign mem_211_6_W0_en = W0_en & W0_addr_sel == 8'hd3;
  assign mem_211_6_W0_mask = W0_mask[6];
  assign mem_211_7_R0_addr = R0_addr[25:0];
  assign mem_211_7_R0_clk = R0_clk;
  assign mem_211_7_R0_en = R0_en & R0_addr_sel == 8'hd3;
  assign mem_211_7_W0_addr = W0_addr[25:0];
  assign mem_211_7_W0_clk = W0_clk;
  assign mem_211_7_W0_data = W0_data[63:56];
  assign mem_211_7_W0_en = W0_en & W0_addr_sel == 8'hd3;
  assign mem_211_7_W0_mask = W0_mask[7];
  assign mem_212_0_R0_addr = R0_addr[25:0];
  assign mem_212_0_R0_clk = R0_clk;
  assign mem_212_0_R0_en = R0_en & R0_addr_sel == 8'hd4;
  assign mem_212_0_W0_addr = W0_addr[25:0];
  assign mem_212_0_W0_clk = W0_clk;
  assign mem_212_0_W0_data = W0_data[7:0];
  assign mem_212_0_W0_en = W0_en & W0_addr_sel == 8'hd4;
  assign mem_212_0_W0_mask = W0_mask[0];
  assign mem_212_1_R0_addr = R0_addr[25:0];
  assign mem_212_1_R0_clk = R0_clk;
  assign mem_212_1_R0_en = R0_en & R0_addr_sel == 8'hd4;
  assign mem_212_1_W0_addr = W0_addr[25:0];
  assign mem_212_1_W0_clk = W0_clk;
  assign mem_212_1_W0_data = W0_data[15:8];
  assign mem_212_1_W0_en = W0_en & W0_addr_sel == 8'hd4;
  assign mem_212_1_W0_mask = W0_mask[1];
  assign mem_212_2_R0_addr = R0_addr[25:0];
  assign mem_212_2_R0_clk = R0_clk;
  assign mem_212_2_R0_en = R0_en & R0_addr_sel == 8'hd4;
  assign mem_212_2_W0_addr = W0_addr[25:0];
  assign mem_212_2_W0_clk = W0_clk;
  assign mem_212_2_W0_data = W0_data[23:16];
  assign mem_212_2_W0_en = W0_en & W0_addr_sel == 8'hd4;
  assign mem_212_2_W0_mask = W0_mask[2];
  assign mem_212_3_R0_addr = R0_addr[25:0];
  assign mem_212_3_R0_clk = R0_clk;
  assign mem_212_3_R0_en = R0_en & R0_addr_sel == 8'hd4;
  assign mem_212_3_W0_addr = W0_addr[25:0];
  assign mem_212_3_W0_clk = W0_clk;
  assign mem_212_3_W0_data = W0_data[31:24];
  assign mem_212_3_W0_en = W0_en & W0_addr_sel == 8'hd4;
  assign mem_212_3_W0_mask = W0_mask[3];
  assign mem_212_4_R0_addr = R0_addr[25:0];
  assign mem_212_4_R0_clk = R0_clk;
  assign mem_212_4_R0_en = R0_en & R0_addr_sel == 8'hd4;
  assign mem_212_4_W0_addr = W0_addr[25:0];
  assign mem_212_4_W0_clk = W0_clk;
  assign mem_212_4_W0_data = W0_data[39:32];
  assign mem_212_4_W0_en = W0_en & W0_addr_sel == 8'hd4;
  assign mem_212_4_W0_mask = W0_mask[4];
  assign mem_212_5_R0_addr = R0_addr[25:0];
  assign mem_212_5_R0_clk = R0_clk;
  assign mem_212_5_R0_en = R0_en & R0_addr_sel == 8'hd4;
  assign mem_212_5_W0_addr = W0_addr[25:0];
  assign mem_212_5_W0_clk = W0_clk;
  assign mem_212_5_W0_data = W0_data[47:40];
  assign mem_212_5_W0_en = W0_en & W0_addr_sel == 8'hd4;
  assign mem_212_5_W0_mask = W0_mask[5];
  assign mem_212_6_R0_addr = R0_addr[25:0];
  assign mem_212_6_R0_clk = R0_clk;
  assign mem_212_6_R0_en = R0_en & R0_addr_sel == 8'hd4;
  assign mem_212_6_W0_addr = W0_addr[25:0];
  assign mem_212_6_W0_clk = W0_clk;
  assign mem_212_6_W0_data = W0_data[55:48];
  assign mem_212_6_W0_en = W0_en & W0_addr_sel == 8'hd4;
  assign mem_212_6_W0_mask = W0_mask[6];
  assign mem_212_7_R0_addr = R0_addr[25:0];
  assign mem_212_7_R0_clk = R0_clk;
  assign mem_212_7_R0_en = R0_en & R0_addr_sel == 8'hd4;
  assign mem_212_7_W0_addr = W0_addr[25:0];
  assign mem_212_7_W0_clk = W0_clk;
  assign mem_212_7_W0_data = W0_data[63:56];
  assign mem_212_7_W0_en = W0_en & W0_addr_sel == 8'hd4;
  assign mem_212_7_W0_mask = W0_mask[7];
  assign mem_213_0_R0_addr = R0_addr[25:0];
  assign mem_213_0_R0_clk = R0_clk;
  assign mem_213_0_R0_en = R0_en & R0_addr_sel == 8'hd5;
  assign mem_213_0_W0_addr = W0_addr[25:0];
  assign mem_213_0_W0_clk = W0_clk;
  assign mem_213_0_W0_data = W0_data[7:0];
  assign mem_213_0_W0_en = W0_en & W0_addr_sel == 8'hd5;
  assign mem_213_0_W0_mask = W0_mask[0];
  assign mem_213_1_R0_addr = R0_addr[25:0];
  assign mem_213_1_R0_clk = R0_clk;
  assign mem_213_1_R0_en = R0_en & R0_addr_sel == 8'hd5;
  assign mem_213_1_W0_addr = W0_addr[25:0];
  assign mem_213_1_W0_clk = W0_clk;
  assign mem_213_1_W0_data = W0_data[15:8];
  assign mem_213_1_W0_en = W0_en & W0_addr_sel == 8'hd5;
  assign mem_213_1_W0_mask = W0_mask[1];
  assign mem_213_2_R0_addr = R0_addr[25:0];
  assign mem_213_2_R0_clk = R0_clk;
  assign mem_213_2_R0_en = R0_en & R0_addr_sel == 8'hd5;
  assign mem_213_2_W0_addr = W0_addr[25:0];
  assign mem_213_2_W0_clk = W0_clk;
  assign mem_213_2_W0_data = W0_data[23:16];
  assign mem_213_2_W0_en = W0_en & W0_addr_sel == 8'hd5;
  assign mem_213_2_W0_mask = W0_mask[2];
  assign mem_213_3_R0_addr = R0_addr[25:0];
  assign mem_213_3_R0_clk = R0_clk;
  assign mem_213_3_R0_en = R0_en & R0_addr_sel == 8'hd5;
  assign mem_213_3_W0_addr = W0_addr[25:0];
  assign mem_213_3_W0_clk = W0_clk;
  assign mem_213_3_W0_data = W0_data[31:24];
  assign mem_213_3_W0_en = W0_en & W0_addr_sel == 8'hd5;
  assign mem_213_3_W0_mask = W0_mask[3];
  assign mem_213_4_R0_addr = R0_addr[25:0];
  assign mem_213_4_R0_clk = R0_clk;
  assign mem_213_4_R0_en = R0_en & R0_addr_sel == 8'hd5;
  assign mem_213_4_W0_addr = W0_addr[25:0];
  assign mem_213_4_W0_clk = W0_clk;
  assign mem_213_4_W0_data = W0_data[39:32];
  assign mem_213_4_W0_en = W0_en & W0_addr_sel == 8'hd5;
  assign mem_213_4_W0_mask = W0_mask[4];
  assign mem_213_5_R0_addr = R0_addr[25:0];
  assign mem_213_5_R0_clk = R0_clk;
  assign mem_213_5_R0_en = R0_en & R0_addr_sel == 8'hd5;
  assign mem_213_5_W0_addr = W0_addr[25:0];
  assign mem_213_5_W0_clk = W0_clk;
  assign mem_213_5_W0_data = W0_data[47:40];
  assign mem_213_5_W0_en = W0_en & W0_addr_sel == 8'hd5;
  assign mem_213_5_W0_mask = W0_mask[5];
  assign mem_213_6_R0_addr = R0_addr[25:0];
  assign mem_213_6_R0_clk = R0_clk;
  assign mem_213_6_R0_en = R0_en & R0_addr_sel == 8'hd5;
  assign mem_213_6_W0_addr = W0_addr[25:0];
  assign mem_213_6_W0_clk = W0_clk;
  assign mem_213_6_W0_data = W0_data[55:48];
  assign mem_213_6_W0_en = W0_en & W0_addr_sel == 8'hd5;
  assign mem_213_6_W0_mask = W0_mask[6];
  assign mem_213_7_R0_addr = R0_addr[25:0];
  assign mem_213_7_R0_clk = R0_clk;
  assign mem_213_7_R0_en = R0_en & R0_addr_sel == 8'hd5;
  assign mem_213_7_W0_addr = W0_addr[25:0];
  assign mem_213_7_W0_clk = W0_clk;
  assign mem_213_7_W0_data = W0_data[63:56];
  assign mem_213_7_W0_en = W0_en & W0_addr_sel == 8'hd5;
  assign mem_213_7_W0_mask = W0_mask[7];
  assign mem_214_0_R0_addr = R0_addr[25:0];
  assign mem_214_0_R0_clk = R0_clk;
  assign mem_214_0_R0_en = R0_en & R0_addr_sel == 8'hd6;
  assign mem_214_0_W0_addr = W0_addr[25:0];
  assign mem_214_0_W0_clk = W0_clk;
  assign mem_214_0_W0_data = W0_data[7:0];
  assign mem_214_0_W0_en = W0_en & W0_addr_sel == 8'hd6;
  assign mem_214_0_W0_mask = W0_mask[0];
  assign mem_214_1_R0_addr = R0_addr[25:0];
  assign mem_214_1_R0_clk = R0_clk;
  assign mem_214_1_R0_en = R0_en & R0_addr_sel == 8'hd6;
  assign mem_214_1_W0_addr = W0_addr[25:0];
  assign mem_214_1_W0_clk = W0_clk;
  assign mem_214_1_W0_data = W0_data[15:8];
  assign mem_214_1_W0_en = W0_en & W0_addr_sel == 8'hd6;
  assign mem_214_1_W0_mask = W0_mask[1];
  assign mem_214_2_R0_addr = R0_addr[25:0];
  assign mem_214_2_R0_clk = R0_clk;
  assign mem_214_2_R0_en = R0_en & R0_addr_sel == 8'hd6;
  assign mem_214_2_W0_addr = W0_addr[25:0];
  assign mem_214_2_W0_clk = W0_clk;
  assign mem_214_2_W0_data = W0_data[23:16];
  assign mem_214_2_W0_en = W0_en & W0_addr_sel == 8'hd6;
  assign mem_214_2_W0_mask = W0_mask[2];
  assign mem_214_3_R0_addr = R0_addr[25:0];
  assign mem_214_3_R0_clk = R0_clk;
  assign mem_214_3_R0_en = R0_en & R0_addr_sel == 8'hd6;
  assign mem_214_3_W0_addr = W0_addr[25:0];
  assign mem_214_3_W0_clk = W0_clk;
  assign mem_214_3_W0_data = W0_data[31:24];
  assign mem_214_3_W0_en = W0_en & W0_addr_sel == 8'hd6;
  assign mem_214_3_W0_mask = W0_mask[3];
  assign mem_214_4_R0_addr = R0_addr[25:0];
  assign mem_214_4_R0_clk = R0_clk;
  assign mem_214_4_R0_en = R0_en & R0_addr_sel == 8'hd6;
  assign mem_214_4_W0_addr = W0_addr[25:0];
  assign mem_214_4_W0_clk = W0_clk;
  assign mem_214_4_W0_data = W0_data[39:32];
  assign mem_214_4_W0_en = W0_en & W0_addr_sel == 8'hd6;
  assign mem_214_4_W0_mask = W0_mask[4];
  assign mem_214_5_R0_addr = R0_addr[25:0];
  assign mem_214_5_R0_clk = R0_clk;
  assign mem_214_5_R0_en = R0_en & R0_addr_sel == 8'hd6;
  assign mem_214_5_W0_addr = W0_addr[25:0];
  assign mem_214_5_W0_clk = W0_clk;
  assign mem_214_5_W0_data = W0_data[47:40];
  assign mem_214_5_W0_en = W0_en & W0_addr_sel == 8'hd6;
  assign mem_214_5_W0_mask = W0_mask[5];
  assign mem_214_6_R0_addr = R0_addr[25:0];
  assign mem_214_6_R0_clk = R0_clk;
  assign mem_214_6_R0_en = R0_en & R0_addr_sel == 8'hd6;
  assign mem_214_6_W0_addr = W0_addr[25:0];
  assign mem_214_6_W0_clk = W0_clk;
  assign mem_214_6_W0_data = W0_data[55:48];
  assign mem_214_6_W0_en = W0_en & W0_addr_sel == 8'hd6;
  assign mem_214_6_W0_mask = W0_mask[6];
  assign mem_214_7_R0_addr = R0_addr[25:0];
  assign mem_214_7_R0_clk = R0_clk;
  assign mem_214_7_R0_en = R0_en & R0_addr_sel == 8'hd6;
  assign mem_214_7_W0_addr = W0_addr[25:0];
  assign mem_214_7_W0_clk = W0_clk;
  assign mem_214_7_W0_data = W0_data[63:56];
  assign mem_214_7_W0_en = W0_en & W0_addr_sel == 8'hd6;
  assign mem_214_7_W0_mask = W0_mask[7];
  assign mem_215_0_R0_addr = R0_addr[25:0];
  assign mem_215_0_R0_clk = R0_clk;
  assign mem_215_0_R0_en = R0_en & R0_addr_sel == 8'hd7;
  assign mem_215_0_W0_addr = W0_addr[25:0];
  assign mem_215_0_W0_clk = W0_clk;
  assign mem_215_0_W0_data = W0_data[7:0];
  assign mem_215_0_W0_en = W0_en & W0_addr_sel == 8'hd7;
  assign mem_215_0_W0_mask = W0_mask[0];
  assign mem_215_1_R0_addr = R0_addr[25:0];
  assign mem_215_1_R0_clk = R0_clk;
  assign mem_215_1_R0_en = R0_en & R0_addr_sel == 8'hd7;
  assign mem_215_1_W0_addr = W0_addr[25:0];
  assign mem_215_1_W0_clk = W0_clk;
  assign mem_215_1_W0_data = W0_data[15:8];
  assign mem_215_1_W0_en = W0_en & W0_addr_sel == 8'hd7;
  assign mem_215_1_W0_mask = W0_mask[1];
  assign mem_215_2_R0_addr = R0_addr[25:0];
  assign mem_215_2_R0_clk = R0_clk;
  assign mem_215_2_R0_en = R0_en & R0_addr_sel == 8'hd7;
  assign mem_215_2_W0_addr = W0_addr[25:0];
  assign mem_215_2_W0_clk = W0_clk;
  assign mem_215_2_W0_data = W0_data[23:16];
  assign mem_215_2_W0_en = W0_en & W0_addr_sel == 8'hd7;
  assign mem_215_2_W0_mask = W0_mask[2];
  assign mem_215_3_R0_addr = R0_addr[25:0];
  assign mem_215_3_R0_clk = R0_clk;
  assign mem_215_3_R0_en = R0_en & R0_addr_sel == 8'hd7;
  assign mem_215_3_W0_addr = W0_addr[25:0];
  assign mem_215_3_W0_clk = W0_clk;
  assign mem_215_3_W0_data = W0_data[31:24];
  assign mem_215_3_W0_en = W0_en & W0_addr_sel == 8'hd7;
  assign mem_215_3_W0_mask = W0_mask[3];
  assign mem_215_4_R0_addr = R0_addr[25:0];
  assign mem_215_4_R0_clk = R0_clk;
  assign mem_215_4_R0_en = R0_en & R0_addr_sel == 8'hd7;
  assign mem_215_4_W0_addr = W0_addr[25:0];
  assign mem_215_4_W0_clk = W0_clk;
  assign mem_215_4_W0_data = W0_data[39:32];
  assign mem_215_4_W0_en = W0_en & W0_addr_sel == 8'hd7;
  assign mem_215_4_W0_mask = W0_mask[4];
  assign mem_215_5_R0_addr = R0_addr[25:0];
  assign mem_215_5_R0_clk = R0_clk;
  assign mem_215_5_R0_en = R0_en & R0_addr_sel == 8'hd7;
  assign mem_215_5_W0_addr = W0_addr[25:0];
  assign mem_215_5_W0_clk = W0_clk;
  assign mem_215_5_W0_data = W0_data[47:40];
  assign mem_215_5_W0_en = W0_en & W0_addr_sel == 8'hd7;
  assign mem_215_5_W0_mask = W0_mask[5];
  assign mem_215_6_R0_addr = R0_addr[25:0];
  assign mem_215_6_R0_clk = R0_clk;
  assign mem_215_6_R0_en = R0_en & R0_addr_sel == 8'hd7;
  assign mem_215_6_W0_addr = W0_addr[25:0];
  assign mem_215_6_W0_clk = W0_clk;
  assign mem_215_6_W0_data = W0_data[55:48];
  assign mem_215_6_W0_en = W0_en & W0_addr_sel == 8'hd7;
  assign mem_215_6_W0_mask = W0_mask[6];
  assign mem_215_7_R0_addr = R0_addr[25:0];
  assign mem_215_7_R0_clk = R0_clk;
  assign mem_215_7_R0_en = R0_en & R0_addr_sel == 8'hd7;
  assign mem_215_7_W0_addr = W0_addr[25:0];
  assign mem_215_7_W0_clk = W0_clk;
  assign mem_215_7_W0_data = W0_data[63:56];
  assign mem_215_7_W0_en = W0_en & W0_addr_sel == 8'hd7;
  assign mem_215_7_W0_mask = W0_mask[7];
  assign mem_216_0_R0_addr = R0_addr[25:0];
  assign mem_216_0_R0_clk = R0_clk;
  assign mem_216_0_R0_en = R0_en & R0_addr_sel == 8'hd8;
  assign mem_216_0_W0_addr = W0_addr[25:0];
  assign mem_216_0_W0_clk = W0_clk;
  assign mem_216_0_W0_data = W0_data[7:0];
  assign mem_216_0_W0_en = W0_en & W0_addr_sel == 8'hd8;
  assign mem_216_0_W0_mask = W0_mask[0];
  assign mem_216_1_R0_addr = R0_addr[25:0];
  assign mem_216_1_R0_clk = R0_clk;
  assign mem_216_1_R0_en = R0_en & R0_addr_sel == 8'hd8;
  assign mem_216_1_W0_addr = W0_addr[25:0];
  assign mem_216_1_W0_clk = W0_clk;
  assign mem_216_1_W0_data = W0_data[15:8];
  assign mem_216_1_W0_en = W0_en & W0_addr_sel == 8'hd8;
  assign mem_216_1_W0_mask = W0_mask[1];
  assign mem_216_2_R0_addr = R0_addr[25:0];
  assign mem_216_2_R0_clk = R0_clk;
  assign mem_216_2_R0_en = R0_en & R0_addr_sel == 8'hd8;
  assign mem_216_2_W0_addr = W0_addr[25:0];
  assign mem_216_2_W0_clk = W0_clk;
  assign mem_216_2_W0_data = W0_data[23:16];
  assign mem_216_2_W0_en = W0_en & W0_addr_sel == 8'hd8;
  assign mem_216_2_W0_mask = W0_mask[2];
  assign mem_216_3_R0_addr = R0_addr[25:0];
  assign mem_216_3_R0_clk = R0_clk;
  assign mem_216_3_R0_en = R0_en & R0_addr_sel == 8'hd8;
  assign mem_216_3_W0_addr = W0_addr[25:0];
  assign mem_216_3_W0_clk = W0_clk;
  assign mem_216_3_W0_data = W0_data[31:24];
  assign mem_216_3_W0_en = W0_en & W0_addr_sel == 8'hd8;
  assign mem_216_3_W0_mask = W0_mask[3];
  assign mem_216_4_R0_addr = R0_addr[25:0];
  assign mem_216_4_R0_clk = R0_clk;
  assign mem_216_4_R0_en = R0_en & R0_addr_sel == 8'hd8;
  assign mem_216_4_W0_addr = W0_addr[25:0];
  assign mem_216_4_W0_clk = W0_clk;
  assign mem_216_4_W0_data = W0_data[39:32];
  assign mem_216_4_W0_en = W0_en & W0_addr_sel == 8'hd8;
  assign mem_216_4_W0_mask = W0_mask[4];
  assign mem_216_5_R0_addr = R0_addr[25:0];
  assign mem_216_5_R0_clk = R0_clk;
  assign mem_216_5_R0_en = R0_en & R0_addr_sel == 8'hd8;
  assign mem_216_5_W0_addr = W0_addr[25:0];
  assign mem_216_5_W0_clk = W0_clk;
  assign mem_216_5_W0_data = W0_data[47:40];
  assign mem_216_5_W0_en = W0_en & W0_addr_sel == 8'hd8;
  assign mem_216_5_W0_mask = W0_mask[5];
  assign mem_216_6_R0_addr = R0_addr[25:0];
  assign mem_216_6_R0_clk = R0_clk;
  assign mem_216_6_R0_en = R0_en & R0_addr_sel == 8'hd8;
  assign mem_216_6_W0_addr = W0_addr[25:0];
  assign mem_216_6_W0_clk = W0_clk;
  assign mem_216_6_W0_data = W0_data[55:48];
  assign mem_216_6_W0_en = W0_en & W0_addr_sel == 8'hd8;
  assign mem_216_6_W0_mask = W0_mask[6];
  assign mem_216_7_R0_addr = R0_addr[25:0];
  assign mem_216_7_R0_clk = R0_clk;
  assign mem_216_7_R0_en = R0_en & R0_addr_sel == 8'hd8;
  assign mem_216_7_W0_addr = W0_addr[25:0];
  assign mem_216_7_W0_clk = W0_clk;
  assign mem_216_7_W0_data = W0_data[63:56];
  assign mem_216_7_W0_en = W0_en & W0_addr_sel == 8'hd8;
  assign mem_216_7_W0_mask = W0_mask[7];
  assign mem_217_0_R0_addr = R0_addr[25:0];
  assign mem_217_0_R0_clk = R0_clk;
  assign mem_217_0_R0_en = R0_en & R0_addr_sel == 8'hd9;
  assign mem_217_0_W0_addr = W0_addr[25:0];
  assign mem_217_0_W0_clk = W0_clk;
  assign mem_217_0_W0_data = W0_data[7:0];
  assign mem_217_0_W0_en = W0_en & W0_addr_sel == 8'hd9;
  assign mem_217_0_W0_mask = W0_mask[0];
  assign mem_217_1_R0_addr = R0_addr[25:0];
  assign mem_217_1_R0_clk = R0_clk;
  assign mem_217_1_R0_en = R0_en & R0_addr_sel == 8'hd9;
  assign mem_217_1_W0_addr = W0_addr[25:0];
  assign mem_217_1_W0_clk = W0_clk;
  assign mem_217_1_W0_data = W0_data[15:8];
  assign mem_217_1_W0_en = W0_en & W0_addr_sel == 8'hd9;
  assign mem_217_1_W0_mask = W0_mask[1];
  assign mem_217_2_R0_addr = R0_addr[25:0];
  assign mem_217_2_R0_clk = R0_clk;
  assign mem_217_2_R0_en = R0_en & R0_addr_sel == 8'hd9;
  assign mem_217_2_W0_addr = W0_addr[25:0];
  assign mem_217_2_W0_clk = W0_clk;
  assign mem_217_2_W0_data = W0_data[23:16];
  assign mem_217_2_W0_en = W0_en & W0_addr_sel == 8'hd9;
  assign mem_217_2_W0_mask = W0_mask[2];
  assign mem_217_3_R0_addr = R0_addr[25:0];
  assign mem_217_3_R0_clk = R0_clk;
  assign mem_217_3_R0_en = R0_en & R0_addr_sel == 8'hd9;
  assign mem_217_3_W0_addr = W0_addr[25:0];
  assign mem_217_3_W0_clk = W0_clk;
  assign mem_217_3_W0_data = W0_data[31:24];
  assign mem_217_3_W0_en = W0_en & W0_addr_sel == 8'hd9;
  assign mem_217_3_W0_mask = W0_mask[3];
  assign mem_217_4_R0_addr = R0_addr[25:0];
  assign mem_217_4_R0_clk = R0_clk;
  assign mem_217_4_R0_en = R0_en & R0_addr_sel == 8'hd9;
  assign mem_217_4_W0_addr = W0_addr[25:0];
  assign mem_217_4_W0_clk = W0_clk;
  assign mem_217_4_W0_data = W0_data[39:32];
  assign mem_217_4_W0_en = W0_en & W0_addr_sel == 8'hd9;
  assign mem_217_4_W0_mask = W0_mask[4];
  assign mem_217_5_R0_addr = R0_addr[25:0];
  assign mem_217_5_R0_clk = R0_clk;
  assign mem_217_5_R0_en = R0_en & R0_addr_sel == 8'hd9;
  assign mem_217_5_W0_addr = W0_addr[25:0];
  assign mem_217_5_W0_clk = W0_clk;
  assign mem_217_5_W0_data = W0_data[47:40];
  assign mem_217_5_W0_en = W0_en & W0_addr_sel == 8'hd9;
  assign mem_217_5_W0_mask = W0_mask[5];
  assign mem_217_6_R0_addr = R0_addr[25:0];
  assign mem_217_6_R0_clk = R0_clk;
  assign mem_217_6_R0_en = R0_en & R0_addr_sel == 8'hd9;
  assign mem_217_6_W0_addr = W0_addr[25:0];
  assign mem_217_6_W0_clk = W0_clk;
  assign mem_217_6_W0_data = W0_data[55:48];
  assign mem_217_6_W0_en = W0_en & W0_addr_sel == 8'hd9;
  assign mem_217_6_W0_mask = W0_mask[6];
  assign mem_217_7_R0_addr = R0_addr[25:0];
  assign mem_217_7_R0_clk = R0_clk;
  assign mem_217_7_R0_en = R0_en & R0_addr_sel == 8'hd9;
  assign mem_217_7_W0_addr = W0_addr[25:0];
  assign mem_217_7_W0_clk = W0_clk;
  assign mem_217_7_W0_data = W0_data[63:56];
  assign mem_217_7_W0_en = W0_en & W0_addr_sel == 8'hd9;
  assign mem_217_7_W0_mask = W0_mask[7];
  assign mem_218_0_R0_addr = R0_addr[25:0];
  assign mem_218_0_R0_clk = R0_clk;
  assign mem_218_0_R0_en = R0_en & R0_addr_sel == 8'hda;
  assign mem_218_0_W0_addr = W0_addr[25:0];
  assign mem_218_0_W0_clk = W0_clk;
  assign mem_218_0_W0_data = W0_data[7:0];
  assign mem_218_0_W0_en = W0_en & W0_addr_sel == 8'hda;
  assign mem_218_0_W0_mask = W0_mask[0];
  assign mem_218_1_R0_addr = R0_addr[25:0];
  assign mem_218_1_R0_clk = R0_clk;
  assign mem_218_1_R0_en = R0_en & R0_addr_sel == 8'hda;
  assign mem_218_1_W0_addr = W0_addr[25:0];
  assign mem_218_1_W0_clk = W0_clk;
  assign mem_218_1_W0_data = W0_data[15:8];
  assign mem_218_1_W0_en = W0_en & W0_addr_sel == 8'hda;
  assign mem_218_1_W0_mask = W0_mask[1];
  assign mem_218_2_R0_addr = R0_addr[25:0];
  assign mem_218_2_R0_clk = R0_clk;
  assign mem_218_2_R0_en = R0_en & R0_addr_sel == 8'hda;
  assign mem_218_2_W0_addr = W0_addr[25:0];
  assign mem_218_2_W0_clk = W0_clk;
  assign mem_218_2_W0_data = W0_data[23:16];
  assign mem_218_2_W0_en = W0_en & W0_addr_sel == 8'hda;
  assign mem_218_2_W0_mask = W0_mask[2];
  assign mem_218_3_R0_addr = R0_addr[25:0];
  assign mem_218_3_R0_clk = R0_clk;
  assign mem_218_3_R0_en = R0_en & R0_addr_sel == 8'hda;
  assign mem_218_3_W0_addr = W0_addr[25:0];
  assign mem_218_3_W0_clk = W0_clk;
  assign mem_218_3_W0_data = W0_data[31:24];
  assign mem_218_3_W0_en = W0_en & W0_addr_sel == 8'hda;
  assign mem_218_3_W0_mask = W0_mask[3];
  assign mem_218_4_R0_addr = R0_addr[25:0];
  assign mem_218_4_R0_clk = R0_clk;
  assign mem_218_4_R0_en = R0_en & R0_addr_sel == 8'hda;
  assign mem_218_4_W0_addr = W0_addr[25:0];
  assign mem_218_4_W0_clk = W0_clk;
  assign mem_218_4_W0_data = W0_data[39:32];
  assign mem_218_4_W0_en = W0_en & W0_addr_sel == 8'hda;
  assign mem_218_4_W0_mask = W0_mask[4];
  assign mem_218_5_R0_addr = R0_addr[25:0];
  assign mem_218_5_R0_clk = R0_clk;
  assign mem_218_5_R0_en = R0_en & R0_addr_sel == 8'hda;
  assign mem_218_5_W0_addr = W0_addr[25:0];
  assign mem_218_5_W0_clk = W0_clk;
  assign mem_218_5_W0_data = W0_data[47:40];
  assign mem_218_5_W0_en = W0_en & W0_addr_sel == 8'hda;
  assign mem_218_5_W0_mask = W0_mask[5];
  assign mem_218_6_R0_addr = R0_addr[25:0];
  assign mem_218_6_R0_clk = R0_clk;
  assign mem_218_6_R0_en = R0_en & R0_addr_sel == 8'hda;
  assign mem_218_6_W0_addr = W0_addr[25:0];
  assign mem_218_6_W0_clk = W0_clk;
  assign mem_218_6_W0_data = W0_data[55:48];
  assign mem_218_6_W0_en = W0_en & W0_addr_sel == 8'hda;
  assign mem_218_6_W0_mask = W0_mask[6];
  assign mem_218_7_R0_addr = R0_addr[25:0];
  assign mem_218_7_R0_clk = R0_clk;
  assign mem_218_7_R0_en = R0_en & R0_addr_sel == 8'hda;
  assign mem_218_7_W0_addr = W0_addr[25:0];
  assign mem_218_7_W0_clk = W0_clk;
  assign mem_218_7_W0_data = W0_data[63:56];
  assign mem_218_7_W0_en = W0_en & W0_addr_sel == 8'hda;
  assign mem_218_7_W0_mask = W0_mask[7];
  assign mem_219_0_R0_addr = R0_addr[25:0];
  assign mem_219_0_R0_clk = R0_clk;
  assign mem_219_0_R0_en = R0_en & R0_addr_sel == 8'hdb;
  assign mem_219_0_W0_addr = W0_addr[25:0];
  assign mem_219_0_W0_clk = W0_clk;
  assign mem_219_0_W0_data = W0_data[7:0];
  assign mem_219_0_W0_en = W0_en & W0_addr_sel == 8'hdb;
  assign mem_219_0_W0_mask = W0_mask[0];
  assign mem_219_1_R0_addr = R0_addr[25:0];
  assign mem_219_1_R0_clk = R0_clk;
  assign mem_219_1_R0_en = R0_en & R0_addr_sel == 8'hdb;
  assign mem_219_1_W0_addr = W0_addr[25:0];
  assign mem_219_1_W0_clk = W0_clk;
  assign mem_219_1_W0_data = W0_data[15:8];
  assign mem_219_1_W0_en = W0_en & W0_addr_sel == 8'hdb;
  assign mem_219_1_W0_mask = W0_mask[1];
  assign mem_219_2_R0_addr = R0_addr[25:0];
  assign mem_219_2_R0_clk = R0_clk;
  assign mem_219_2_R0_en = R0_en & R0_addr_sel == 8'hdb;
  assign mem_219_2_W0_addr = W0_addr[25:0];
  assign mem_219_2_W0_clk = W0_clk;
  assign mem_219_2_W0_data = W0_data[23:16];
  assign mem_219_2_W0_en = W0_en & W0_addr_sel == 8'hdb;
  assign mem_219_2_W0_mask = W0_mask[2];
  assign mem_219_3_R0_addr = R0_addr[25:0];
  assign mem_219_3_R0_clk = R0_clk;
  assign mem_219_3_R0_en = R0_en & R0_addr_sel == 8'hdb;
  assign mem_219_3_W0_addr = W0_addr[25:0];
  assign mem_219_3_W0_clk = W0_clk;
  assign mem_219_3_W0_data = W0_data[31:24];
  assign mem_219_3_W0_en = W0_en & W0_addr_sel == 8'hdb;
  assign mem_219_3_W0_mask = W0_mask[3];
  assign mem_219_4_R0_addr = R0_addr[25:0];
  assign mem_219_4_R0_clk = R0_clk;
  assign mem_219_4_R0_en = R0_en & R0_addr_sel == 8'hdb;
  assign mem_219_4_W0_addr = W0_addr[25:0];
  assign mem_219_4_W0_clk = W0_clk;
  assign mem_219_4_W0_data = W0_data[39:32];
  assign mem_219_4_W0_en = W0_en & W0_addr_sel == 8'hdb;
  assign mem_219_4_W0_mask = W0_mask[4];
  assign mem_219_5_R0_addr = R0_addr[25:0];
  assign mem_219_5_R0_clk = R0_clk;
  assign mem_219_5_R0_en = R0_en & R0_addr_sel == 8'hdb;
  assign mem_219_5_W0_addr = W0_addr[25:0];
  assign mem_219_5_W0_clk = W0_clk;
  assign mem_219_5_W0_data = W0_data[47:40];
  assign mem_219_5_W0_en = W0_en & W0_addr_sel == 8'hdb;
  assign mem_219_5_W0_mask = W0_mask[5];
  assign mem_219_6_R0_addr = R0_addr[25:0];
  assign mem_219_6_R0_clk = R0_clk;
  assign mem_219_6_R0_en = R0_en & R0_addr_sel == 8'hdb;
  assign mem_219_6_W0_addr = W0_addr[25:0];
  assign mem_219_6_W0_clk = W0_clk;
  assign mem_219_6_W0_data = W0_data[55:48];
  assign mem_219_6_W0_en = W0_en & W0_addr_sel == 8'hdb;
  assign mem_219_6_W0_mask = W0_mask[6];
  assign mem_219_7_R0_addr = R0_addr[25:0];
  assign mem_219_7_R0_clk = R0_clk;
  assign mem_219_7_R0_en = R0_en & R0_addr_sel == 8'hdb;
  assign mem_219_7_W0_addr = W0_addr[25:0];
  assign mem_219_7_W0_clk = W0_clk;
  assign mem_219_7_W0_data = W0_data[63:56];
  assign mem_219_7_W0_en = W0_en & W0_addr_sel == 8'hdb;
  assign mem_219_7_W0_mask = W0_mask[7];
  assign mem_220_0_R0_addr = R0_addr[25:0];
  assign mem_220_0_R0_clk = R0_clk;
  assign mem_220_0_R0_en = R0_en & R0_addr_sel == 8'hdc;
  assign mem_220_0_W0_addr = W0_addr[25:0];
  assign mem_220_0_W0_clk = W0_clk;
  assign mem_220_0_W0_data = W0_data[7:0];
  assign mem_220_0_W0_en = W0_en & W0_addr_sel == 8'hdc;
  assign mem_220_0_W0_mask = W0_mask[0];
  assign mem_220_1_R0_addr = R0_addr[25:0];
  assign mem_220_1_R0_clk = R0_clk;
  assign mem_220_1_R0_en = R0_en & R0_addr_sel == 8'hdc;
  assign mem_220_1_W0_addr = W0_addr[25:0];
  assign mem_220_1_W0_clk = W0_clk;
  assign mem_220_1_W0_data = W0_data[15:8];
  assign mem_220_1_W0_en = W0_en & W0_addr_sel == 8'hdc;
  assign mem_220_1_W0_mask = W0_mask[1];
  assign mem_220_2_R0_addr = R0_addr[25:0];
  assign mem_220_2_R0_clk = R0_clk;
  assign mem_220_2_R0_en = R0_en & R0_addr_sel == 8'hdc;
  assign mem_220_2_W0_addr = W0_addr[25:0];
  assign mem_220_2_W0_clk = W0_clk;
  assign mem_220_2_W0_data = W0_data[23:16];
  assign mem_220_2_W0_en = W0_en & W0_addr_sel == 8'hdc;
  assign mem_220_2_W0_mask = W0_mask[2];
  assign mem_220_3_R0_addr = R0_addr[25:0];
  assign mem_220_3_R0_clk = R0_clk;
  assign mem_220_3_R0_en = R0_en & R0_addr_sel == 8'hdc;
  assign mem_220_3_W0_addr = W0_addr[25:0];
  assign mem_220_3_W0_clk = W0_clk;
  assign mem_220_3_W0_data = W0_data[31:24];
  assign mem_220_3_W0_en = W0_en & W0_addr_sel == 8'hdc;
  assign mem_220_3_W0_mask = W0_mask[3];
  assign mem_220_4_R0_addr = R0_addr[25:0];
  assign mem_220_4_R0_clk = R0_clk;
  assign mem_220_4_R0_en = R0_en & R0_addr_sel == 8'hdc;
  assign mem_220_4_W0_addr = W0_addr[25:0];
  assign mem_220_4_W0_clk = W0_clk;
  assign mem_220_4_W0_data = W0_data[39:32];
  assign mem_220_4_W0_en = W0_en & W0_addr_sel == 8'hdc;
  assign mem_220_4_W0_mask = W0_mask[4];
  assign mem_220_5_R0_addr = R0_addr[25:0];
  assign mem_220_5_R0_clk = R0_clk;
  assign mem_220_5_R0_en = R0_en & R0_addr_sel == 8'hdc;
  assign mem_220_5_W0_addr = W0_addr[25:0];
  assign mem_220_5_W0_clk = W0_clk;
  assign mem_220_5_W0_data = W0_data[47:40];
  assign mem_220_5_W0_en = W0_en & W0_addr_sel == 8'hdc;
  assign mem_220_5_W0_mask = W0_mask[5];
  assign mem_220_6_R0_addr = R0_addr[25:0];
  assign mem_220_6_R0_clk = R0_clk;
  assign mem_220_6_R0_en = R0_en & R0_addr_sel == 8'hdc;
  assign mem_220_6_W0_addr = W0_addr[25:0];
  assign mem_220_6_W0_clk = W0_clk;
  assign mem_220_6_W0_data = W0_data[55:48];
  assign mem_220_6_W0_en = W0_en & W0_addr_sel == 8'hdc;
  assign mem_220_6_W0_mask = W0_mask[6];
  assign mem_220_7_R0_addr = R0_addr[25:0];
  assign mem_220_7_R0_clk = R0_clk;
  assign mem_220_7_R0_en = R0_en & R0_addr_sel == 8'hdc;
  assign mem_220_7_W0_addr = W0_addr[25:0];
  assign mem_220_7_W0_clk = W0_clk;
  assign mem_220_7_W0_data = W0_data[63:56];
  assign mem_220_7_W0_en = W0_en & W0_addr_sel == 8'hdc;
  assign mem_220_7_W0_mask = W0_mask[7];
  assign mem_221_0_R0_addr = R0_addr[25:0];
  assign mem_221_0_R0_clk = R0_clk;
  assign mem_221_0_R0_en = R0_en & R0_addr_sel == 8'hdd;
  assign mem_221_0_W0_addr = W0_addr[25:0];
  assign mem_221_0_W0_clk = W0_clk;
  assign mem_221_0_W0_data = W0_data[7:0];
  assign mem_221_0_W0_en = W0_en & W0_addr_sel == 8'hdd;
  assign mem_221_0_W0_mask = W0_mask[0];
  assign mem_221_1_R0_addr = R0_addr[25:0];
  assign mem_221_1_R0_clk = R0_clk;
  assign mem_221_1_R0_en = R0_en & R0_addr_sel == 8'hdd;
  assign mem_221_1_W0_addr = W0_addr[25:0];
  assign mem_221_1_W0_clk = W0_clk;
  assign mem_221_1_W0_data = W0_data[15:8];
  assign mem_221_1_W0_en = W0_en & W0_addr_sel == 8'hdd;
  assign mem_221_1_W0_mask = W0_mask[1];
  assign mem_221_2_R0_addr = R0_addr[25:0];
  assign mem_221_2_R0_clk = R0_clk;
  assign mem_221_2_R0_en = R0_en & R0_addr_sel == 8'hdd;
  assign mem_221_2_W0_addr = W0_addr[25:0];
  assign mem_221_2_W0_clk = W0_clk;
  assign mem_221_2_W0_data = W0_data[23:16];
  assign mem_221_2_W0_en = W0_en & W0_addr_sel == 8'hdd;
  assign mem_221_2_W0_mask = W0_mask[2];
  assign mem_221_3_R0_addr = R0_addr[25:0];
  assign mem_221_3_R0_clk = R0_clk;
  assign mem_221_3_R0_en = R0_en & R0_addr_sel == 8'hdd;
  assign mem_221_3_W0_addr = W0_addr[25:0];
  assign mem_221_3_W0_clk = W0_clk;
  assign mem_221_3_W0_data = W0_data[31:24];
  assign mem_221_3_W0_en = W0_en & W0_addr_sel == 8'hdd;
  assign mem_221_3_W0_mask = W0_mask[3];
  assign mem_221_4_R0_addr = R0_addr[25:0];
  assign mem_221_4_R0_clk = R0_clk;
  assign mem_221_4_R0_en = R0_en & R0_addr_sel == 8'hdd;
  assign mem_221_4_W0_addr = W0_addr[25:0];
  assign mem_221_4_W0_clk = W0_clk;
  assign mem_221_4_W0_data = W0_data[39:32];
  assign mem_221_4_W0_en = W0_en & W0_addr_sel == 8'hdd;
  assign mem_221_4_W0_mask = W0_mask[4];
  assign mem_221_5_R0_addr = R0_addr[25:0];
  assign mem_221_5_R0_clk = R0_clk;
  assign mem_221_5_R0_en = R0_en & R0_addr_sel == 8'hdd;
  assign mem_221_5_W0_addr = W0_addr[25:0];
  assign mem_221_5_W0_clk = W0_clk;
  assign mem_221_5_W0_data = W0_data[47:40];
  assign mem_221_5_W0_en = W0_en & W0_addr_sel == 8'hdd;
  assign mem_221_5_W0_mask = W0_mask[5];
  assign mem_221_6_R0_addr = R0_addr[25:0];
  assign mem_221_6_R0_clk = R0_clk;
  assign mem_221_6_R0_en = R0_en & R0_addr_sel == 8'hdd;
  assign mem_221_6_W0_addr = W0_addr[25:0];
  assign mem_221_6_W0_clk = W0_clk;
  assign mem_221_6_W0_data = W0_data[55:48];
  assign mem_221_6_W0_en = W0_en & W0_addr_sel == 8'hdd;
  assign mem_221_6_W0_mask = W0_mask[6];
  assign mem_221_7_R0_addr = R0_addr[25:0];
  assign mem_221_7_R0_clk = R0_clk;
  assign mem_221_7_R0_en = R0_en & R0_addr_sel == 8'hdd;
  assign mem_221_7_W0_addr = W0_addr[25:0];
  assign mem_221_7_W0_clk = W0_clk;
  assign mem_221_7_W0_data = W0_data[63:56];
  assign mem_221_7_W0_en = W0_en & W0_addr_sel == 8'hdd;
  assign mem_221_7_W0_mask = W0_mask[7];
  assign mem_222_0_R0_addr = R0_addr[25:0];
  assign mem_222_0_R0_clk = R0_clk;
  assign mem_222_0_R0_en = R0_en & R0_addr_sel == 8'hde;
  assign mem_222_0_W0_addr = W0_addr[25:0];
  assign mem_222_0_W0_clk = W0_clk;
  assign mem_222_0_W0_data = W0_data[7:0];
  assign mem_222_0_W0_en = W0_en & W0_addr_sel == 8'hde;
  assign mem_222_0_W0_mask = W0_mask[0];
  assign mem_222_1_R0_addr = R0_addr[25:0];
  assign mem_222_1_R0_clk = R0_clk;
  assign mem_222_1_R0_en = R0_en & R0_addr_sel == 8'hde;
  assign mem_222_1_W0_addr = W0_addr[25:0];
  assign mem_222_1_W0_clk = W0_clk;
  assign mem_222_1_W0_data = W0_data[15:8];
  assign mem_222_1_W0_en = W0_en & W0_addr_sel == 8'hde;
  assign mem_222_1_W0_mask = W0_mask[1];
  assign mem_222_2_R0_addr = R0_addr[25:0];
  assign mem_222_2_R0_clk = R0_clk;
  assign mem_222_2_R0_en = R0_en & R0_addr_sel == 8'hde;
  assign mem_222_2_W0_addr = W0_addr[25:0];
  assign mem_222_2_W0_clk = W0_clk;
  assign mem_222_2_W0_data = W0_data[23:16];
  assign mem_222_2_W0_en = W0_en & W0_addr_sel == 8'hde;
  assign mem_222_2_W0_mask = W0_mask[2];
  assign mem_222_3_R0_addr = R0_addr[25:0];
  assign mem_222_3_R0_clk = R0_clk;
  assign mem_222_3_R0_en = R0_en & R0_addr_sel == 8'hde;
  assign mem_222_3_W0_addr = W0_addr[25:0];
  assign mem_222_3_W0_clk = W0_clk;
  assign mem_222_3_W0_data = W0_data[31:24];
  assign mem_222_3_W0_en = W0_en & W0_addr_sel == 8'hde;
  assign mem_222_3_W0_mask = W0_mask[3];
  assign mem_222_4_R0_addr = R0_addr[25:0];
  assign mem_222_4_R0_clk = R0_clk;
  assign mem_222_4_R0_en = R0_en & R0_addr_sel == 8'hde;
  assign mem_222_4_W0_addr = W0_addr[25:0];
  assign mem_222_4_W0_clk = W0_clk;
  assign mem_222_4_W0_data = W0_data[39:32];
  assign mem_222_4_W0_en = W0_en & W0_addr_sel == 8'hde;
  assign mem_222_4_W0_mask = W0_mask[4];
  assign mem_222_5_R0_addr = R0_addr[25:0];
  assign mem_222_5_R0_clk = R0_clk;
  assign mem_222_5_R0_en = R0_en & R0_addr_sel == 8'hde;
  assign mem_222_5_W0_addr = W0_addr[25:0];
  assign mem_222_5_W0_clk = W0_clk;
  assign mem_222_5_W0_data = W0_data[47:40];
  assign mem_222_5_W0_en = W0_en & W0_addr_sel == 8'hde;
  assign mem_222_5_W0_mask = W0_mask[5];
  assign mem_222_6_R0_addr = R0_addr[25:0];
  assign mem_222_6_R0_clk = R0_clk;
  assign mem_222_6_R0_en = R0_en & R0_addr_sel == 8'hde;
  assign mem_222_6_W0_addr = W0_addr[25:0];
  assign mem_222_6_W0_clk = W0_clk;
  assign mem_222_6_W0_data = W0_data[55:48];
  assign mem_222_6_W0_en = W0_en & W0_addr_sel == 8'hde;
  assign mem_222_6_W0_mask = W0_mask[6];
  assign mem_222_7_R0_addr = R0_addr[25:0];
  assign mem_222_7_R0_clk = R0_clk;
  assign mem_222_7_R0_en = R0_en & R0_addr_sel == 8'hde;
  assign mem_222_7_W0_addr = W0_addr[25:0];
  assign mem_222_7_W0_clk = W0_clk;
  assign mem_222_7_W0_data = W0_data[63:56];
  assign mem_222_7_W0_en = W0_en & W0_addr_sel == 8'hde;
  assign mem_222_7_W0_mask = W0_mask[7];
  assign mem_223_0_R0_addr = R0_addr[25:0];
  assign mem_223_0_R0_clk = R0_clk;
  assign mem_223_0_R0_en = R0_en & R0_addr_sel == 8'hdf;
  assign mem_223_0_W0_addr = W0_addr[25:0];
  assign mem_223_0_W0_clk = W0_clk;
  assign mem_223_0_W0_data = W0_data[7:0];
  assign mem_223_0_W0_en = W0_en & W0_addr_sel == 8'hdf;
  assign mem_223_0_W0_mask = W0_mask[0];
  assign mem_223_1_R0_addr = R0_addr[25:0];
  assign mem_223_1_R0_clk = R0_clk;
  assign mem_223_1_R0_en = R0_en & R0_addr_sel == 8'hdf;
  assign mem_223_1_W0_addr = W0_addr[25:0];
  assign mem_223_1_W0_clk = W0_clk;
  assign mem_223_1_W0_data = W0_data[15:8];
  assign mem_223_1_W0_en = W0_en & W0_addr_sel == 8'hdf;
  assign mem_223_1_W0_mask = W0_mask[1];
  assign mem_223_2_R0_addr = R0_addr[25:0];
  assign mem_223_2_R0_clk = R0_clk;
  assign mem_223_2_R0_en = R0_en & R0_addr_sel == 8'hdf;
  assign mem_223_2_W0_addr = W0_addr[25:0];
  assign mem_223_2_W0_clk = W0_clk;
  assign mem_223_2_W0_data = W0_data[23:16];
  assign mem_223_2_W0_en = W0_en & W0_addr_sel == 8'hdf;
  assign mem_223_2_W0_mask = W0_mask[2];
  assign mem_223_3_R0_addr = R0_addr[25:0];
  assign mem_223_3_R0_clk = R0_clk;
  assign mem_223_3_R0_en = R0_en & R0_addr_sel == 8'hdf;
  assign mem_223_3_W0_addr = W0_addr[25:0];
  assign mem_223_3_W0_clk = W0_clk;
  assign mem_223_3_W0_data = W0_data[31:24];
  assign mem_223_3_W0_en = W0_en & W0_addr_sel == 8'hdf;
  assign mem_223_3_W0_mask = W0_mask[3];
  assign mem_223_4_R0_addr = R0_addr[25:0];
  assign mem_223_4_R0_clk = R0_clk;
  assign mem_223_4_R0_en = R0_en & R0_addr_sel == 8'hdf;
  assign mem_223_4_W0_addr = W0_addr[25:0];
  assign mem_223_4_W0_clk = W0_clk;
  assign mem_223_4_W0_data = W0_data[39:32];
  assign mem_223_4_W0_en = W0_en & W0_addr_sel == 8'hdf;
  assign mem_223_4_W0_mask = W0_mask[4];
  assign mem_223_5_R0_addr = R0_addr[25:0];
  assign mem_223_5_R0_clk = R0_clk;
  assign mem_223_5_R0_en = R0_en & R0_addr_sel == 8'hdf;
  assign mem_223_5_W0_addr = W0_addr[25:0];
  assign mem_223_5_W0_clk = W0_clk;
  assign mem_223_5_W0_data = W0_data[47:40];
  assign mem_223_5_W0_en = W0_en & W0_addr_sel == 8'hdf;
  assign mem_223_5_W0_mask = W0_mask[5];
  assign mem_223_6_R0_addr = R0_addr[25:0];
  assign mem_223_6_R0_clk = R0_clk;
  assign mem_223_6_R0_en = R0_en & R0_addr_sel == 8'hdf;
  assign mem_223_6_W0_addr = W0_addr[25:0];
  assign mem_223_6_W0_clk = W0_clk;
  assign mem_223_6_W0_data = W0_data[55:48];
  assign mem_223_6_W0_en = W0_en & W0_addr_sel == 8'hdf;
  assign mem_223_6_W0_mask = W0_mask[6];
  assign mem_223_7_R0_addr = R0_addr[25:0];
  assign mem_223_7_R0_clk = R0_clk;
  assign mem_223_7_R0_en = R0_en & R0_addr_sel == 8'hdf;
  assign mem_223_7_W0_addr = W0_addr[25:0];
  assign mem_223_7_W0_clk = W0_clk;
  assign mem_223_7_W0_data = W0_data[63:56];
  assign mem_223_7_W0_en = W0_en & W0_addr_sel == 8'hdf;
  assign mem_223_7_W0_mask = W0_mask[7];
  assign mem_224_0_R0_addr = R0_addr[25:0];
  assign mem_224_0_R0_clk = R0_clk;
  assign mem_224_0_R0_en = R0_en & R0_addr_sel == 8'he0;
  assign mem_224_0_W0_addr = W0_addr[25:0];
  assign mem_224_0_W0_clk = W0_clk;
  assign mem_224_0_W0_data = W0_data[7:0];
  assign mem_224_0_W0_en = W0_en & W0_addr_sel == 8'he0;
  assign mem_224_0_W0_mask = W0_mask[0];
  assign mem_224_1_R0_addr = R0_addr[25:0];
  assign mem_224_1_R0_clk = R0_clk;
  assign mem_224_1_R0_en = R0_en & R0_addr_sel == 8'he0;
  assign mem_224_1_W0_addr = W0_addr[25:0];
  assign mem_224_1_W0_clk = W0_clk;
  assign mem_224_1_W0_data = W0_data[15:8];
  assign mem_224_1_W0_en = W0_en & W0_addr_sel == 8'he0;
  assign mem_224_1_W0_mask = W0_mask[1];
  assign mem_224_2_R0_addr = R0_addr[25:0];
  assign mem_224_2_R0_clk = R0_clk;
  assign mem_224_2_R0_en = R0_en & R0_addr_sel == 8'he0;
  assign mem_224_2_W0_addr = W0_addr[25:0];
  assign mem_224_2_W0_clk = W0_clk;
  assign mem_224_2_W0_data = W0_data[23:16];
  assign mem_224_2_W0_en = W0_en & W0_addr_sel == 8'he0;
  assign mem_224_2_W0_mask = W0_mask[2];
  assign mem_224_3_R0_addr = R0_addr[25:0];
  assign mem_224_3_R0_clk = R0_clk;
  assign mem_224_3_R0_en = R0_en & R0_addr_sel == 8'he0;
  assign mem_224_3_W0_addr = W0_addr[25:0];
  assign mem_224_3_W0_clk = W0_clk;
  assign mem_224_3_W0_data = W0_data[31:24];
  assign mem_224_3_W0_en = W0_en & W0_addr_sel == 8'he0;
  assign mem_224_3_W0_mask = W0_mask[3];
  assign mem_224_4_R0_addr = R0_addr[25:0];
  assign mem_224_4_R0_clk = R0_clk;
  assign mem_224_4_R0_en = R0_en & R0_addr_sel == 8'he0;
  assign mem_224_4_W0_addr = W0_addr[25:0];
  assign mem_224_4_W0_clk = W0_clk;
  assign mem_224_4_W0_data = W0_data[39:32];
  assign mem_224_4_W0_en = W0_en & W0_addr_sel == 8'he0;
  assign mem_224_4_W0_mask = W0_mask[4];
  assign mem_224_5_R0_addr = R0_addr[25:0];
  assign mem_224_5_R0_clk = R0_clk;
  assign mem_224_5_R0_en = R0_en & R0_addr_sel == 8'he0;
  assign mem_224_5_W0_addr = W0_addr[25:0];
  assign mem_224_5_W0_clk = W0_clk;
  assign mem_224_5_W0_data = W0_data[47:40];
  assign mem_224_5_W0_en = W0_en & W0_addr_sel == 8'he0;
  assign mem_224_5_W0_mask = W0_mask[5];
  assign mem_224_6_R0_addr = R0_addr[25:0];
  assign mem_224_6_R0_clk = R0_clk;
  assign mem_224_6_R0_en = R0_en & R0_addr_sel == 8'he0;
  assign mem_224_6_W0_addr = W0_addr[25:0];
  assign mem_224_6_W0_clk = W0_clk;
  assign mem_224_6_W0_data = W0_data[55:48];
  assign mem_224_6_W0_en = W0_en & W0_addr_sel == 8'he0;
  assign mem_224_6_W0_mask = W0_mask[6];
  assign mem_224_7_R0_addr = R0_addr[25:0];
  assign mem_224_7_R0_clk = R0_clk;
  assign mem_224_7_R0_en = R0_en & R0_addr_sel == 8'he0;
  assign mem_224_7_W0_addr = W0_addr[25:0];
  assign mem_224_7_W0_clk = W0_clk;
  assign mem_224_7_W0_data = W0_data[63:56];
  assign mem_224_7_W0_en = W0_en & W0_addr_sel == 8'he0;
  assign mem_224_7_W0_mask = W0_mask[7];
  assign mem_225_0_R0_addr = R0_addr[25:0];
  assign mem_225_0_R0_clk = R0_clk;
  assign mem_225_0_R0_en = R0_en & R0_addr_sel == 8'he1;
  assign mem_225_0_W0_addr = W0_addr[25:0];
  assign mem_225_0_W0_clk = W0_clk;
  assign mem_225_0_W0_data = W0_data[7:0];
  assign mem_225_0_W0_en = W0_en & W0_addr_sel == 8'he1;
  assign mem_225_0_W0_mask = W0_mask[0];
  assign mem_225_1_R0_addr = R0_addr[25:0];
  assign mem_225_1_R0_clk = R0_clk;
  assign mem_225_1_R0_en = R0_en & R0_addr_sel == 8'he1;
  assign mem_225_1_W0_addr = W0_addr[25:0];
  assign mem_225_1_W0_clk = W0_clk;
  assign mem_225_1_W0_data = W0_data[15:8];
  assign mem_225_1_W0_en = W0_en & W0_addr_sel == 8'he1;
  assign mem_225_1_W0_mask = W0_mask[1];
  assign mem_225_2_R0_addr = R0_addr[25:0];
  assign mem_225_2_R0_clk = R0_clk;
  assign mem_225_2_R0_en = R0_en & R0_addr_sel == 8'he1;
  assign mem_225_2_W0_addr = W0_addr[25:0];
  assign mem_225_2_W0_clk = W0_clk;
  assign mem_225_2_W0_data = W0_data[23:16];
  assign mem_225_2_W0_en = W0_en & W0_addr_sel == 8'he1;
  assign mem_225_2_W0_mask = W0_mask[2];
  assign mem_225_3_R0_addr = R0_addr[25:0];
  assign mem_225_3_R0_clk = R0_clk;
  assign mem_225_3_R0_en = R0_en & R0_addr_sel == 8'he1;
  assign mem_225_3_W0_addr = W0_addr[25:0];
  assign mem_225_3_W0_clk = W0_clk;
  assign mem_225_3_W0_data = W0_data[31:24];
  assign mem_225_3_W0_en = W0_en & W0_addr_sel == 8'he1;
  assign mem_225_3_W0_mask = W0_mask[3];
  assign mem_225_4_R0_addr = R0_addr[25:0];
  assign mem_225_4_R0_clk = R0_clk;
  assign mem_225_4_R0_en = R0_en & R0_addr_sel == 8'he1;
  assign mem_225_4_W0_addr = W0_addr[25:0];
  assign mem_225_4_W0_clk = W0_clk;
  assign mem_225_4_W0_data = W0_data[39:32];
  assign mem_225_4_W0_en = W0_en & W0_addr_sel == 8'he1;
  assign mem_225_4_W0_mask = W0_mask[4];
  assign mem_225_5_R0_addr = R0_addr[25:0];
  assign mem_225_5_R0_clk = R0_clk;
  assign mem_225_5_R0_en = R0_en & R0_addr_sel == 8'he1;
  assign mem_225_5_W0_addr = W0_addr[25:0];
  assign mem_225_5_W0_clk = W0_clk;
  assign mem_225_5_W0_data = W0_data[47:40];
  assign mem_225_5_W0_en = W0_en & W0_addr_sel == 8'he1;
  assign mem_225_5_W0_mask = W0_mask[5];
  assign mem_225_6_R0_addr = R0_addr[25:0];
  assign mem_225_6_R0_clk = R0_clk;
  assign mem_225_6_R0_en = R0_en & R0_addr_sel == 8'he1;
  assign mem_225_6_W0_addr = W0_addr[25:0];
  assign mem_225_6_W0_clk = W0_clk;
  assign mem_225_6_W0_data = W0_data[55:48];
  assign mem_225_6_W0_en = W0_en & W0_addr_sel == 8'he1;
  assign mem_225_6_W0_mask = W0_mask[6];
  assign mem_225_7_R0_addr = R0_addr[25:0];
  assign mem_225_7_R0_clk = R0_clk;
  assign mem_225_7_R0_en = R0_en & R0_addr_sel == 8'he1;
  assign mem_225_7_W0_addr = W0_addr[25:0];
  assign mem_225_7_W0_clk = W0_clk;
  assign mem_225_7_W0_data = W0_data[63:56];
  assign mem_225_7_W0_en = W0_en & W0_addr_sel == 8'he1;
  assign mem_225_7_W0_mask = W0_mask[7];
  assign mem_226_0_R0_addr = R0_addr[25:0];
  assign mem_226_0_R0_clk = R0_clk;
  assign mem_226_0_R0_en = R0_en & R0_addr_sel == 8'he2;
  assign mem_226_0_W0_addr = W0_addr[25:0];
  assign mem_226_0_W0_clk = W0_clk;
  assign mem_226_0_W0_data = W0_data[7:0];
  assign mem_226_0_W0_en = W0_en & W0_addr_sel == 8'he2;
  assign mem_226_0_W0_mask = W0_mask[0];
  assign mem_226_1_R0_addr = R0_addr[25:0];
  assign mem_226_1_R0_clk = R0_clk;
  assign mem_226_1_R0_en = R0_en & R0_addr_sel == 8'he2;
  assign mem_226_1_W0_addr = W0_addr[25:0];
  assign mem_226_1_W0_clk = W0_clk;
  assign mem_226_1_W0_data = W0_data[15:8];
  assign mem_226_1_W0_en = W0_en & W0_addr_sel == 8'he2;
  assign mem_226_1_W0_mask = W0_mask[1];
  assign mem_226_2_R0_addr = R0_addr[25:0];
  assign mem_226_2_R0_clk = R0_clk;
  assign mem_226_2_R0_en = R0_en & R0_addr_sel == 8'he2;
  assign mem_226_2_W0_addr = W0_addr[25:0];
  assign mem_226_2_W0_clk = W0_clk;
  assign mem_226_2_W0_data = W0_data[23:16];
  assign mem_226_2_W0_en = W0_en & W0_addr_sel == 8'he2;
  assign mem_226_2_W0_mask = W0_mask[2];
  assign mem_226_3_R0_addr = R0_addr[25:0];
  assign mem_226_3_R0_clk = R0_clk;
  assign mem_226_3_R0_en = R0_en & R0_addr_sel == 8'he2;
  assign mem_226_3_W0_addr = W0_addr[25:0];
  assign mem_226_3_W0_clk = W0_clk;
  assign mem_226_3_W0_data = W0_data[31:24];
  assign mem_226_3_W0_en = W0_en & W0_addr_sel == 8'he2;
  assign mem_226_3_W0_mask = W0_mask[3];
  assign mem_226_4_R0_addr = R0_addr[25:0];
  assign mem_226_4_R0_clk = R0_clk;
  assign mem_226_4_R0_en = R0_en & R0_addr_sel == 8'he2;
  assign mem_226_4_W0_addr = W0_addr[25:0];
  assign mem_226_4_W0_clk = W0_clk;
  assign mem_226_4_W0_data = W0_data[39:32];
  assign mem_226_4_W0_en = W0_en & W0_addr_sel == 8'he2;
  assign mem_226_4_W0_mask = W0_mask[4];
  assign mem_226_5_R0_addr = R0_addr[25:0];
  assign mem_226_5_R0_clk = R0_clk;
  assign mem_226_5_R0_en = R0_en & R0_addr_sel == 8'he2;
  assign mem_226_5_W0_addr = W0_addr[25:0];
  assign mem_226_5_W0_clk = W0_clk;
  assign mem_226_5_W0_data = W0_data[47:40];
  assign mem_226_5_W0_en = W0_en & W0_addr_sel == 8'he2;
  assign mem_226_5_W0_mask = W0_mask[5];
  assign mem_226_6_R0_addr = R0_addr[25:0];
  assign mem_226_6_R0_clk = R0_clk;
  assign mem_226_6_R0_en = R0_en & R0_addr_sel == 8'he2;
  assign mem_226_6_W0_addr = W0_addr[25:0];
  assign mem_226_6_W0_clk = W0_clk;
  assign mem_226_6_W0_data = W0_data[55:48];
  assign mem_226_6_W0_en = W0_en & W0_addr_sel == 8'he2;
  assign mem_226_6_W0_mask = W0_mask[6];
  assign mem_226_7_R0_addr = R0_addr[25:0];
  assign mem_226_7_R0_clk = R0_clk;
  assign mem_226_7_R0_en = R0_en & R0_addr_sel == 8'he2;
  assign mem_226_7_W0_addr = W0_addr[25:0];
  assign mem_226_7_W0_clk = W0_clk;
  assign mem_226_7_W0_data = W0_data[63:56];
  assign mem_226_7_W0_en = W0_en & W0_addr_sel == 8'he2;
  assign mem_226_7_W0_mask = W0_mask[7];
  assign mem_227_0_R0_addr = R0_addr[25:0];
  assign mem_227_0_R0_clk = R0_clk;
  assign mem_227_0_R0_en = R0_en & R0_addr_sel == 8'he3;
  assign mem_227_0_W0_addr = W0_addr[25:0];
  assign mem_227_0_W0_clk = W0_clk;
  assign mem_227_0_W0_data = W0_data[7:0];
  assign mem_227_0_W0_en = W0_en & W0_addr_sel == 8'he3;
  assign mem_227_0_W0_mask = W0_mask[0];
  assign mem_227_1_R0_addr = R0_addr[25:0];
  assign mem_227_1_R0_clk = R0_clk;
  assign mem_227_1_R0_en = R0_en & R0_addr_sel == 8'he3;
  assign mem_227_1_W0_addr = W0_addr[25:0];
  assign mem_227_1_W0_clk = W0_clk;
  assign mem_227_1_W0_data = W0_data[15:8];
  assign mem_227_1_W0_en = W0_en & W0_addr_sel == 8'he3;
  assign mem_227_1_W0_mask = W0_mask[1];
  assign mem_227_2_R0_addr = R0_addr[25:0];
  assign mem_227_2_R0_clk = R0_clk;
  assign mem_227_2_R0_en = R0_en & R0_addr_sel == 8'he3;
  assign mem_227_2_W0_addr = W0_addr[25:0];
  assign mem_227_2_W0_clk = W0_clk;
  assign mem_227_2_W0_data = W0_data[23:16];
  assign mem_227_2_W0_en = W0_en & W0_addr_sel == 8'he3;
  assign mem_227_2_W0_mask = W0_mask[2];
  assign mem_227_3_R0_addr = R0_addr[25:0];
  assign mem_227_3_R0_clk = R0_clk;
  assign mem_227_3_R0_en = R0_en & R0_addr_sel == 8'he3;
  assign mem_227_3_W0_addr = W0_addr[25:0];
  assign mem_227_3_W0_clk = W0_clk;
  assign mem_227_3_W0_data = W0_data[31:24];
  assign mem_227_3_W0_en = W0_en & W0_addr_sel == 8'he3;
  assign mem_227_3_W0_mask = W0_mask[3];
  assign mem_227_4_R0_addr = R0_addr[25:0];
  assign mem_227_4_R0_clk = R0_clk;
  assign mem_227_4_R0_en = R0_en & R0_addr_sel == 8'he3;
  assign mem_227_4_W0_addr = W0_addr[25:0];
  assign mem_227_4_W0_clk = W0_clk;
  assign mem_227_4_W0_data = W0_data[39:32];
  assign mem_227_4_W0_en = W0_en & W0_addr_sel == 8'he3;
  assign mem_227_4_W0_mask = W0_mask[4];
  assign mem_227_5_R0_addr = R0_addr[25:0];
  assign mem_227_5_R0_clk = R0_clk;
  assign mem_227_5_R0_en = R0_en & R0_addr_sel == 8'he3;
  assign mem_227_5_W0_addr = W0_addr[25:0];
  assign mem_227_5_W0_clk = W0_clk;
  assign mem_227_5_W0_data = W0_data[47:40];
  assign mem_227_5_W0_en = W0_en & W0_addr_sel == 8'he3;
  assign mem_227_5_W0_mask = W0_mask[5];
  assign mem_227_6_R0_addr = R0_addr[25:0];
  assign mem_227_6_R0_clk = R0_clk;
  assign mem_227_6_R0_en = R0_en & R0_addr_sel == 8'he3;
  assign mem_227_6_W0_addr = W0_addr[25:0];
  assign mem_227_6_W0_clk = W0_clk;
  assign mem_227_6_W0_data = W0_data[55:48];
  assign mem_227_6_W0_en = W0_en & W0_addr_sel == 8'he3;
  assign mem_227_6_W0_mask = W0_mask[6];
  assign mem_227_7_R0_addr = R0_addr[25:0];
  assign mem_227_7_R0_clk = R0_clk;
  assign mem_227_7_R0_en = R0_en & R0_addr_sel == 8'he3;
  assign mem_227_7_W0_addr = W0_addr[25:0];
  assign mem_227_7_W0_clk = W0_clk;
  assign mem_227_7_W0_data = W0_data[63:56];
  assign mem_227_7_W0_en = W0_en & W0_addr_sel == 8'he3;
  assign mem_227_7_W0_mask = W0_mask[7];
  assign mem_228_0_R0_addr = R0_addr[25:0];
  assign mem_228_0_R0_clk = R0_clk;
  assign mem_228_0_R0_en = R0_en & R0_addr_sel == 8'he4;
  assign mem_228_0_W0_addr = W0_addr[25:0];
  assign mem_228_0_W0_clk = W0_clk;
  assign mem_228_0_W0_data = W0_data[7:0];
  assign mem_228_0_W0_en = W0_en & W0_addr_sel == 8'he4;
  assign mem_228_0_W0_mask = W0_mask[0];
  assign mem_228_1_R0_addr = R0_addr[25:0];
  assign mem_228_1_R0_clk = R0_clk;
  assign mem_228_1_R0_en = R0_en & R0_addr_sel == 8'he4;
  assign mem_228_1_W0_addr = W0_addr[25:0];
  assign mem_228_1_W0_clk = W0_clk;
  assign mem_228_1_W0_data = W0_data[15:8];
  assign mem_228_1_W0_en = W0_en & W0_addr_sel == 8'he4;
  assign mem_228_1_W0_mask = W0_mask[1];
  assign mem_228_2_R0_addr = R0_addr[25:0];
  assign mem_228_2_R0_clk = R0_clk;
  assign mem_228_2_R0_en = R0_en & R0_addr_sel == 8'he4;
  assign mem_228_2_W0_addr = W0_addr[25:0];
  assign mem_228_2_W0_clk = W0_clk;
  assign mem_228_2_W0_data = W0_data[23:16];
  assign mem_228_2_W0_en = W0_en & W0_addr_sel == 8'he4;
  assign mem_228_2_W0_mask = W0_mask[2];
  assign mem_228_3_R0_addr = R0_addr[25:0];
  assign mem_228_3_R0_clk = R0_clk;
  assign mem_228_3_R0_en = R0_en & R0_addr_sel == 8'he4;
  assign mem_228_3_W0_addr = W0_addr[25:0];
  assign mem_228_3_W0_clk = W0_clk;
  assign mem_228_3_W0_data = W0_data[31:24];
  assign mem_228_3_W0_en = W0_en & W0_addr_sel == 8'he4;
  assign mem_228_3_W0_mask = W0_mask[3];
  assign mem_228_4_R0_addr = R0_addr[25:0];
  assign mem_228_4_R0_clk = R0_clk;
  assign mem_228_4_R0_en = R0_en & R0_addr_sel == 8'he4;
  assign mem_228_4_W0_addr = W0_addr[25:0];
  assign mem_228_4_W0_clk = W0_clk;
  assign mem_228_4_W0_data = W0_data[39:32];
  assign mem_228_4_W0_en = W0_en & W0_addr_sel == 8'he4;
  assign mem_228_4_W0_mask = W0_mask[4];
  assign mem_228_5_R0_addr = R0_addr[25:0];
  assign mem_228_5_R0_clk = R0_clk;
  assign mem_228_5_R0_en = R0_en & R0_addr_sel == 8'he4;
  assign mem_228_5_W0_addr = W0_addr[25:0];
  assign mem_228_5_W0_clk = W0_clk;
  assign mem_228_5_W0_data = W0_data[47:40];
  assign mem_228_5_W0_en = W0_en & W0_addr_sel == 8'he4;
  assign mem_228_5_W0_mask = W0_mask[5];
  assign mem_228_6_R0_addr = R0_addr[25:0];
  assign mem_228_6_R0_clk = R0_clk;
  assign mem_228_6_R0_en = R0_en & R0_addr_sel == 8'he4;
  assign mem_228_6_W0_addr = W0_addr[25:0];
  assign mem_228_6_W0_clk = W0_clk;
  assign mem_228_6_W0_data = W0_data[55:48];
  assign mem_228_6_W0_en = W0_en & W0_addr_sel == 8'he4;
  assign mem_228_6_W0_mask = W0_mask[6];
  assign mem_228_7_R0_addr = R0_addr[25:0];
  assign mem_228_7_R0_clk = R0_clk;
  assign mem_228_7_R0_en = R0_en & R0_addr_sel == 8'he4;
  assign mem_228_7_W0_addr = W0_addr[25:0];
  assign mem_228_7_W0_clk = W0_clk;
  assign mem_228_7_W0_data = W0_data[63:56];
  assign mem_228_7_W0_en = W0_en & W0_addr_sel == 8'he4;
  assign mem_228_7_W0_mask = W0_mask[7];
  assign mem_229_0_R0_addr = R0_addr[25:0];
  assign mem_229_0_R0_clk = R0_clk;
  assign mem_229_0_R0_en = R0_en & R0_addr_sel == 8'he5;
  assign mem_229_0_W0_addr = W0_addr[25:0];
  assign mem_229_0_W0_clk = W0_clk;
  assign mem_229_0_W0_data = W0_data[7:0];
  assign mem_229_0_W0_en = W0_en & W0_addr_sel == 8'he5;
  assign mem_229_0_W0_mask = W0_mask[0];
  assign mem_229_1_R0_addr = R0_addr[25:0];
  assign mem_229_1_R0_clk = R0_clk;
  assign mem_229_1_R0_en = R0_en & R0_addr_sel == 8'he5;
  assign mem_229_1_W0_addr = W0_addr[25:0];
  assign mem_229_1_W0_clk = W0_clk;
  assign mem_229_1_W0_data = W0_data[15:8];
  assign mem_229_1_W0_en = W0_en & W0_addr_sel == 8'he5;
  assign mem_229_1_W0_mask = W0_mask[1];
  assign mem_229_2_R0_addr = R0_addr[25:0];
  assign mem_229_2_R0_clk = R0_clk;
  assign mem_229_2_R0_en = R0_en & R0_addr_sel == 8'he5;
  assign mem_229_2_W0_addr = W0_addr[25:0];
  assign mem_229_2_W0_clk = W0_clk;
  assign mem_229_2_W0_data = W0_data[23:16];
  assign mem_229_2_W0_en = W0_en & W0_addr_sel == 8'he5;
  assign mem_229_2_W0_mask = W0_mask[2];
  assign mem_229_3_R0_addr = R0_addr[25:0];
  assign mem_229_3_R0_clk = R0_clk;
  assign mem_229_3_R0_en = R0_en & R0_addr_sel == 8'he5;
  assign mem_229_3_W0_addr = W0_addr[25:0];
  assign mem_229_3_W0_clk = W0_clk;
  assign mem_229_3_W0_data = W0_data[31:24];
  assign mem_229_3_W0_en = W0_en & W0_addr_sel == 8'he5;
  assign mem_229_3_W0_mask = W0_mask[3];
  assign mem_229_4_R0_addr = R0_addr[25:0];
  assign mem_229_4_R0_clk = R0_clk;
  assign mem_229_4_R0_en = R0_en & R0_addr_sel == 8'he5;
  assign mem_229_4_W0_addr = W0_addr[25:0];
  assign mem_229_4_W0_clk = W0_clk;
  assign mem_229_4_W0_data = W0_data[39:32];
  assign mem_229_4_W0_en = W0_en & W0_addr_sel == 8'he5;
  assign mem_229_4_W0_mask = W0_mask[4];
  assign mem_229_5_R0_addr = R0_addr[25:0];
  assign mem_229_5_R0_clk = R0_clk;
  assign mem_229_5_R0_en = R0_en & R0_addr_sel == 8'he5;
  assign mem_229_5_W0_addr = W0_addr[25:0];
  assign mem_229_5_W0_clk = W0_clk;
  assign mem_229_5_W0_data = W0_data[47:40];
  assign mem_229_5_W0_en = W0_en & W0_addr_sel == 8'he5;
  assign mem_229_5_W0_mask = W0_mask[5];
  assign mem_229_6_R0_addr = R0_addr[25:0];
  assign mem_229_6_R0_clk = R0_clk;
  assign mem_229_6_R0_en = R0_en & R0_addr_sel == 8'he5;
  assign mem_229_6_W0_addr = W0_addr[25:0];
  assign mem_229_6_W0_clk = W0_clk;
  assign mem_229_6_W0_data = W0_data[55:48];
  assign mem_229_6_W0_en = W0_en & W0_addr_sel == 8'he5;
  assign mem_229_6_W0_mask = W0_mask[6];
  assign mem_229_7_R0_addr = R0_addr[25:0];
  assign mem_229_7_R0_clk = R0_clk;
  assign mem_229_7_R0_en = R0_en & R0_addr_sel == 8'he5;
  assign mem_229_7_W0_addr = W0_addr[25:0];
  assign mem_229_7_W0_clk = W0_clk;
  assign mem_229_7_W0_data = W0_data[63:56];
  assign mem_229_7_W0_en = W0_en & W0_addr_sel == 8'he5;
  assign mem_229_7_W0_mask = W0_mask[7];
  assign mem_230_0_R0_addr = R0_addr[25:0];
  assign mem_230_0_R0_clk = R0_clk;
  assign mem_230_0_R0_en = R0_en & R0_addr_sel == 8'he6;
  assign mem_230_0_W0_addr = W0_addr[25:0];
  assign mem_230_0_W0_clk = W0_clk;
  assign mem_230_0_W0_data = W0_data[7:0];
  assign mem_230_0_W0_en = W0_en & W0_addr_sel == 8'he6;
  assign mem_230_0_W0_mask = W0_mask[0];
  assign mem_230_1_R0_addr = R0_addr[25:0];
  assign mem_230_1_R0_clk = R0_clk;
  assign mem_230_1_R0_en = R0_en & R0_addr_sel == 8'he6;
  assign mem_230_1_W0_addr = W0_addr[25:0];
  assign mem_230_1_W0_clk = W0_clk;
  assign mem_230_1_W0_data = W0_data[15:8];
  assign mem_230_1_W0_en = W0_en & W0_addr_sel == 8'he6;
  assign mem_230_1_W0_mask = W0_mask[1];
  assign mem_230_2_R0_addr = R0_addr[25:0];
  assign mem_230_2_R0_clk = R0_clk;
  assign mem_230_2_R0_en = R0_en & R0_addr_sel == 8'he6;
  assign mem_230_2_W0_addr = W0_addr[25:0];
  assign mem_230_2_W0_clk = W0_clk;
  assign mem_230_2_W0_data = W0_data[23:16];
  assign mem_230_2_W0_en = W0_en & W0_addr_sel == 8'he6;
  assign mem_230_2_W0_mask = W0_mask[2];
  assign mem_230_3_R0_addr = R0_addr[25:0];
  assign mem_230_3_R0_clk = R0_clk;
  assign mem_230_3_R0_en = R0_en & R0_addr_sel == 8'he6;
  assign mem_230_3_W0_addr = W0_addr[25:0];
  assign mem_230_3_W0_clk = W0_clk;
  assign mem_230_3_W0_data = W0_data[31:24];
  assign mem_230_3_W0_en = W0_en & W0_addr_sel == 8'he6;
  assign mem_230_3_W0_mask = W0_mask[3];
  assign mem_230_4_R0_addr = R0_addr[25:0];
  assign mem_230_4_R0_clk = R0_clk;
  assign mem_230_4_R0_en = R0_en & R0_addr_sel == 8'he6;
  assign mem_230_4_W0_addr = W0_addr[25:0];
  assign mem_230_4_W0_clk = W0_clk;
  assign mem_230_4_W0_data = W0_data[39:32];
  assign mem_230_4_W0_en = W0_en & W0_addr_sel == 8'he6;
  assign mem_230_4_W0_mask = W0_mask[4];
  assign mem_230_5_R0_addr = R0_addr[25:0];
  assign mem_230_5_R0_clk = R0_clk;
  assign mem_230_5_R0_en = R0_en & R0_addr_sel == 8'he6;
  assign mem_230_5_W0_addr = W0_addr[25:0];
  assign mem_230_5_W0_clk = W0_clk;
  assign mem_230_5_W0_data = W0_data[47:40];
  assign mem_230_5_W0_en = W0_en & W0_addr_sel == 8'he6;
  assign mem_230_5_W0_mask = W0_mask[5];
  assign mem_230_6_R0_addr = R0_addr[25:0];
  assign mem_230_6_R0_clk = R0_clk;
  assign mem_230_6_R0_en = R0_en & R0_addr_sel == 8'he6;
  assign mem_230_6_W0_addr = W0_addr[25:0];
  assign mem_230_6_W0_clk = W0_clk;
  assign mem_230_6_W0_data = W0_data[55:48];
  assign mem_230_6_W0_en = W0_en & W0_addr_sel == 8'he6;
  assign mem_230_6_W0_mask = W0_mask[6];
  assign mem_230_7_R0_addr = R0_addr[25:0];
  assign mem_230_7_R0_clk = R0_clk;
  assign mem_230_7_R0_en = R0_en & R0_addr_sel == 8'he6;
  assign mem_230_7_W0_addr = W0_addr[25:0];
  assign mem_230_7_W0_clk = W0_clk;
  assign mem_230_7_W0_data = W0_data[63:56];
  assign mem_230_7_W0_en = W0_en & W0_addr_sel == 8'he6;
  assign mem_230_7_W0_mask = W0_mask[7];
  assign mem_231_0_R0_addr = R0_addr[25:0];
  assign mem_231_0_R0_clk = R0_clk;
  assign mem_231_0_R0_en = R0_en & R0_addr_sel == 8'he7;
  assign mem_231_0_W0_addr = W0_addr[25:0];
  assign mem_231_0_W0_clk = W0_clk;
  assign mem_231_0_W0_data = W0_data[7:0];
  assign mem_231_0_W0_en = W0_en & W0_addr_sel == 8'he7;
  assign mem_231_0_W0_mask = W0_mask[0];
  assign mem_231_1_R0_addr = R0_addr[25:0];
  assign mem_231_1_R0_clk = R0_clk;
  assign mem_231_1_R0_en = R0_en & R0_addr_sel == 8'he7;
  assign mem_231_1_W0_addr = W0_addr[25:0];
  assign mem_231_1_W0_clk = W0_clk;
  assign mem_231_1_W0_data = W0_data[15:8];
  assign mem_231_1_W0_en = W0_en & W0_addr_sel == 8'he7;
  assign mem_231_1_W0_mask = W0_mask[1];
  assign mem_231_2_R0_addr = R0_addr[25:0];
  assign mem_231_2_R0_clk = R0_clk;
  assign mem_231_2_R0_en = R0_en & R0_addr_sel == 8'he7;
  assign mem_231_2_W0_addr = W0_addr[25:0];
  assign mem_231_2_W0_clk = W0_clk;
  assign mem_231_2_W0_data = W0_data[23:16];
  assign mem_231_2_W0_en = W0_en & W0_addr_sel == 8'he7;
  assign mem_231_2_W0_mask = W0_mask[2];
  assign mem_231_3_R0_addr = R0_addr[25:0];
  assign mem_231_3_R0_clk = R0_clk;
  assign mem_231_3_R0_en = R0_en & R0_addr_sel == 8'he7;
  assign mem_231_3_W0_addr = W0_addr[25:0];
  assign mem_231_3_W0_clk = W0_clk;
  assign mem_231_3_W0_data = W0_data[31:24];
  assign mem_231_3_W0_en = W0_en & W0_addr_sel == 8'he7;
  assign mem_231_3_W0_mask = W0_mask[3];
  assign mem_231_4_R0_addr = R0_addr[25:0];
  assign mem_231_4_R0_clk = R0_clk;
  assign mem_231_4_R0_en = R0_en & R0_addr_sel == 8'he7;
  assign mem_231_4_W0_addr = W0_addr[25:0];
  assign mem_231_4_W0_clk = W0_clk;
  assign mem_231_4_W0_data = W0_data[39:32];
  assign mem_231_4_W0_en = W0_en & W0_addr_sel == 8'he7;
  assign mem_231_4_W0_mask = W0_mask[4];
  assign mem_231_5_R0_addr = R0_addr[25:0];
  assign mem_231_5_R0_clk = R0_clk;
  assign mem_231_5_R0_en = R0_en & R0_addr_sel == 8'he7;
  assign mem_231_5_W0_addr = W0_addr[25:0];
  assign mem_231_5_W0_clk = W0_clk;
  assign mem_231_5_W0_data = W0_data[47:40];
  assign mem_231_5_W0_en = W0_en & W0_addr_sel == 8'he7;
  assign mem_231_5_W0_mask = W0_mask[5];
  assign mem_231_6_R0_addr = R0_addr[25:0];
  assign mem_231_6_R0_clk = R0_clk;
  assign mem_231_6_R0_en = R0_en & R0_addr_sel == 8'he7;
  assign mem_231_6_W0_addr = W0_addr[25:0];
  assign mem_231_6_W0_clk = W0_clk;
  assign mem_231_6_W0_data = W0_data[55:48];
  assign mem_231_6_W0_en = W0_en & W0_addr_sel == 8'he7;
  assign mem_231_6_W0_mask = W0_mask[6];
  assign mem_231_7_R0_addr = R0_addr[25:0];
  assign mem_231_7_R0_clk = R0_clk;
  assign mem_231_7_R0_en = R0_en & R0_addr_sel == 8'he7;
  assign mem_231_7_W0_addr = W0_addr[25:0];
  assign mem_231_7_W0_clk = W0_clk;
  assign mem_231_7_W0_data = W0_data[63:56];
  assign mem_231_7_W0_en = W0_en & W0_addr_sel == 8'he7;
  assign mem_231_7_W0_mask = W0_mask[7];
  assign mem_232_0_R0_addr = R0_addr[25:0];
  assign mem_232_0_R0_clk = R0_clk;
  assign mem_232_0_R0_en = R0_en & R0_addr_sel == 8'he8;
  assign mem_232_0_W0_addr = W0_addr[25:0];
  assign mem_232_0_W0_clk = W0_clk;
  assign mem_232_0_W0_data = W0_data[7:0];
  assign mem_232_0_W0_en = W0_en & W0_addr_sel == 8'he8;
  assign mem_232_0_W0_mask = W0_mask[0];
  assign mem_232_1_R0_addr = R0_addr[25:0];
  assign mem_232_1_R0_clk = R0_clk;
  assign mem_232_1_R0_en = R0_en & R0_addr_sel == 8'he8;
  assign mem_232_1_W0_addr = W0_addr[25:0];
  assign mem_232_1_W0_clk = W0_clk;
  assign mem_232_1_W0_data = W0_data[15:8];
  assign mem_232_1_W0_en = W0_en & W0_addr_sel == 8'he8;
  assign mem_232_1_W0_mask = W0_mask[1];
  assign mem_232_2_R0_addr = R0_addr[25:0];
  assign mem_232_2_R0_clk = R0_clk;
  assign mem_232_2_R0_en = R0_en & R0_addr_sel == 8'he8;
  assign mem_232_2_W0_addr = W0_addr[25:0];
  assign mem_232_2_W0_clk = W0_clk;
  assign mem_232_2_W0_data = W0_data[23:16];
  assign mem_232_2_W0_en = W0_en & W0_addr_sel == 8'he8;
  assign mem_232_2_W0_mask = W0_mask[2];
  assign mem_232_3_R0_addr = R0_addr[25:0];
  assign mem_232_3_R0_clk = R0_clk;
  assign mem_232_3_R0_en = R0_en & R0_addr_sel == 8'he8;
  assign mem_232_3_W0_addr = W0_addr[25:0];
  assign mem_232_3_W0_clk = W0_clk;
  assign mem_232_3_W0_data = W0_data[31:24];
  assign mem_232_3_W0_en = W0_en & W0_addr_sel == 8'he8;
  assign mem_232_3_W0_mask = W0_mask[3];
  assign mem_232_4_R0_addr = R0_addr[25:0];
  assign mem_232_4_R0_clk = R0_clk;
  assign mem_232_4_R0_en = R0_en & R0_addr_sel == 8'he8;
  assign mem_232_4_W0_addr = W0_addr[25:0];
  assign mem_232_4_W0_clk = W0_clk;
  assign mem_232_4_W0_data = W0_data[39:32];
  assign mem_232_4_W0_en = W0_en & W0_addr_sel == 8'he8;
  assign mem_232_4_W0_mask = W0_mask[4];
  assign mem_232_5_R0_addr = R0_addr[25:0];
  assign mem_232_5_R0_clk = R0_clk;
  assign mem_232_5_R0_en = R0_en & R0_addr_sel == 8'he8;
  assign mem_232_5_W0_addr = W0_addr[25:0];
  assign mem_232_5_W0_clk = W0_clk;
  assign mem_232_5_W0_data = W0_data[47:40];
  assign mem_232_5_W0_en = W0_en & W0_addr_sel == 8'he8;
  assign mem_232_5_W0_mask = W0_mask[5];
  assign mem_232_6_R0_addr = R0_addr[25:0];
  assign mem_232_6_R0_clk = R0_clk;
  assign mem_232_6_R0_en = R0_en & R0_addr_sel == 8'he8;
  assign mem_232_6_W0_addr = W0_addr[25:0];
  assign mem_232_6_W0_clk = W0_clk;
  assign mem_232_6_W0_data = W0_data[55:48];
  assign mem_232_6_W0_en = W0_en & W0_addr_sel == 8'he8;
  assign mem_232_6_W0_mask = W0_mask[6];
  assign mem_232_7_R0_addr = R0_addr[25:0];
  assign mem_232_7_R0_clk = R0_clk;
  assign mem_232_7_R0_en = R0_en & R0_addr_sel == 8'he8;
  assign mem_232_7_W0_addr = W0_addr[25:0];
  assign mem_232_7_W0_clk = W0_clk;
  assign mem_232_7_W0_data = W0_data[63:56];
  assign mem_232_7_W0_en = W0_en & W0_addr_sel == 8'he8;
  assign mem_232_7_W0_mask = W0_mask[7];
  assign mem_233_0_R0_addr = R0_addr[25:0];
  assign mem_233_0_R0_clk = R0_clk;
  assign mem_233_0_R0_en = R0_en & R0_addr_sel == 8'he9;
  assign mem_233_0_W0_addr = W0_addr[25:0];
  assign mem_233_0_W0_clk = W0_clk;
  assign mem_233_0_W0_data = W0_data[7:0];
  assign mem_233_0_W0_en = W0_en & W0_addr_sel == 8'he9;
  assign mem_233_0_W0_mask = W0_mask[0];
  assign mem_233_1_R0_addr = R0_addr[25:0];
  assign mem_233_1_R0_clk = R0_clk;
  assign mem_233_1_R0_en = R0_en & R0_addr_sel == 8'he9;
  assign mem_233_1_W0_addr = W0_addr[25:0];
  assign mem_233_1_W0_clk = W0_clk;
  assign mem_233_1_W0_data = W0_data[15:8];
  assign mem_233_1_W0_en = W0_en & W0_addr_sel == 8'he9;
  assign mem_233_1_W0_mask = W0_mask[1];
  assign mem_233_2_R0_addr = R0_addr[25:0];
  assign mem_233_2_R0_clk = R0_clk;
  assign mem_233_2_R0_en = R0_en & R0_addr_sel == 8'he9;
  assign mem_233_2_W0_addr = W0_addr[25:0];
  assign mem_233_2_W0_clk = W0_clk;
  assign mem_233_2_W0_data = W0_data[23:16];
  assign mem_233_2_W0_en = W0_en & W0_addr_sel == 8'he9;
  assign mem_233_2_W0_mask = W0_mask[2];
  assign mem_233_3_R0_addr = R0_addr[25:0];
  assign mem_233_3_R0_clk = R0_clk;
  assign mem_233_3_R0_en = R0_en & R0_addr_sel == 8'he9;
  assign mem_233_3_W0_addr = W0_addr[25:0];
  assign mem_233_3_W0_clk = W0_clk;
  assign mem_233_3_W0_data = W0_data[31:24];
  assign mem_233_3_W0_en = W0_en & W0_addr_sel == 8'he9;
  assign mem_233_3_W0_mask = W0_mask[3];
  assign mem_233_4_R0_addr = R0_addr[25:0];
  assign mem_233_4_R0_clk = R0_clk;
  assign mem_233_4_R0_en = R0_en & R0_addr_sel == 8'he9;
  assign mem_233_4_W0_addr = W0_addr[25:0];
  assign mem_233_4_W0_clk = W0_clk;
  assign mem_233_4_W0_data = W0_data[39:32];
  assign mem_233_4_W0_en = W0_en & W0_addr_sel == 8'he9;
  assign mem_233_4_W0_mask = W0_mask[4];
  assign mem_233_5_R0_addr = R0_addr[25:0];
  assign mem_233_5_R0_clk = R0_clk;
  assign mem_233_5_R0_en = R0_en & R0_addr_sel == 8'he9;
  assign mem_233_5_W0_addr = W0_addr[25:0];
  assign mem_233_5_W0_clk = W0_clk;
  assign mem_233_5_W0_data = W0_data[47:40];
  assign mem_233_5_W0_en = W0_en & W0_addr_sel == 8'he9;
  assign mem_233_5_W0_mask = W0_mask[5];
  assign mem_233_6_R0_addr = R0_addr[25:0];
  assign mem_233_6_R0_clk = R0_clk;
  assign mem_233_6_R0_en = R0_en & R0_addr_sel == 8'he9;
  assign mem_233_6_W0_addr = W0_addr[25:0];
  assign mem_233_6_W0_clk = W0_clk;
  assign mem_233_6_W0_data = W0_data[55:48];
  assign mem_233_6_W0_en = W0_en & W0_addr_sel == 8'he9;
  assign mem_233_6_W0_mask = W0_mask[6];
  assign mem_233_7_R0_addr = R0_addr[25:0];
  assign mem_233_7_R0_clk = R0_clk;
  assign mem_233_7_R0_en = R0_en & R0_addr_sel == 8'he9;
  assign mem_233_7_W0_addr = W0_addr[25:0];
  assign mem_233_7_W0_clk = W0_clk;
  assign mem_233_7_W0_data = W0_data[63:56];
  assign mem_233_7_W0_en = W0_en & W0_addr_sel == 8'he9;
  assign mem_233_7_W0_mask = W0_mask[7];
  assign mem_234_0_R0_addr = R0_addr[25:0];
  assign mem_234_0_R0_clk = R0_clk;
  assign mem_234_0_R0_en = R0_en & R0_addr_sel == 8'hea;
  assign mem_234_0_W0_addr = W0_addr[25:0];
  assign mem_234_0_W0_clk = W0_clk;
  assign mem_234_0_W0_data = W0_data[7:0];
  assign mem_234_0_W0_en = W0_en & W0_addr_sel == 8'hea;
  assign mem_234_0_W0_mask = W0_mask[0];
  assign mem_234_1_R0_addr = R0_addr[25:0];
  assign mem_234_1_R0_clk = R0_clk;
  assign mem_234_1_R0_en = R0_en & R0_addr_sel == 8'hea;
  assign mem_234_1_W0_addr = W0_addr[25:0];
  assign mem_234_1_W0_clk = W0_clk;
  assign mem_234_1_W0_data = W0_data[15:8];
  assign mem_234_1_W0_en = W0_en & W0_addr_sel == 8'hea;
  assign mem_234_1_W0_mask = W0_mask[1];
  assign mem_234_2_R0_addr = R0_addr[25:0];
  assign mem_234_2_R0_clk = R0_clk;
  assign mem_234_2_R0_en = R0_en & R0_addr_sel == 8'hea;
  assign mem_234_2_W0_addr = W0_addr[25:0];
  assign mem_234_2_W0_clk = W0_clk;
  assign mem_234_2_W0_data = W0_data[23:16];
  assign mem_234_2_W0_en = W0_en & W0_addr_sel == 8'hea;
  assign mem_234_2_W0_mask = W0_mask[2];
  assign mem_234_3_R0_addr = R0_addr[25:0];
  assign mem_234_3_R0_clk = R0_clk;
  assign mem_234_3_R0_en = R0_en & R0_addr_sel == 8'hea;
  assign mem_234_3_W0_addr = W0_addr[25:0];
  assign mem_234_3_W0_clk = W0_clk;
  assign mem_234_3_W0_data = W0_data[31:24];
  assign mem_234_3_W0_en = W0_en & W0_addr_sel == 8'hea;
  assign mem_234_3_W0_mask = W0_mask[3];
  assign mem_234_4_R0_addr = R0_addr[25:0];
  assign mem_234_4_R0_clk = R0_clk;
  assign mem_234_4_R0_en = R0_en & R0_addr_sel == 8'hea;
  assign mem_234_4_W0_addr = W0_addr[25:0];
  assign mem_234_4_W0_clk = W0_clk;
  assign mem_234_4_W0_data = W0_data[39:32];
  assign mem_234_4_W0_en = W0_en & W0_addr_sel == 8'hea;
  assign mem_234_4_W0_mask = W0_mask[4];
  assign mem_234_5_R0_addr = R0_addr[25:0];
  assign mem_234_5_R0_clk = R0_clk;
  assign mem_234_5_R0_en = R0_en & R0_addr_sel == 8'hea;
  assign mem_234_5_W0_addr = W0_addr[25:0];
  assign mem_234_5_W0_clk = W0_clk;
  assign mem_234_5_W0_data = W0_data[47:40];
  assign mem_234_5_W0_en = W0_en & W0_addr_sel == 8'hea;
  assign mem_234_5_W0_mask = W0_mask[5];
  assign mem_234_6_R0_addr = R0_addr[25:0];
  assign mem_234_6_R0_clk = R0_clk;
  assign mem_234_6_R0_en = R0_en & R0_addr_sel == 8'hea;
  assign mem_234_6_W0_addr = W0_addr[25:0];
  assign mem_234_6_W0_clk = W0_clk;
  assign mem_234_6_W0_data = W0_data[55:48];
  assign mem_234_6_W0_en = W0_en & W0_addr_sel == 8'hea;
  assign mem_234_6_W0_mask = W0_mask[6];
  assign mem_234_7_R0_addr = R0_addr[25:0];
  assign mem_234_7_R0_clk = R0_clk;
  assign mem_234_7_R0_en = R0_en & R0_addr_sel == 8'hea;
  assign mem_234_7_W0_addr = W0_addr[25:0];
  assign mem_234_7_W0_clk = W0_clk;
  assign mem_234_7_W0_data = W0_data[63:56];
  assign mem_234_7_W0_en = W0_en & W0_addr_sel == 8'hea;
  assign mem_234_7_W0_mask = W0_mask[7];
  assign mem_235_0_R0_addr = R0_addr[25:0];
  assign mem_235_0_R0_clk = R0_clk;
  assign mem_235_0_R0_en = R0_en & R0_addr_sel == 8'heb;
  assign mem_235_0_W0_addr = W0_addr[25:0];
  assign mem_235_0_W0_clk = W0_clk;
  assign mem_235_0_W0_data = W0_data[7:0];
  assign mem_235_0_W0_en = W0_en & W0_addr_sel == 8'heb;
  assign mem_235_0_W0_mask = W0_mask[0];
  assign mem_235_1_R0_addr = R0_addr[25:0];
  assign mem_235_1_R0_clk = R0_clk;
  assign mem_235_1_R0_en = R0_en & R0_addr_sel == 8'heb;
  assign mem_235_1_W0_addr = W0_addr[25:0];
  assign mem_235_1_W0_clk = W0_clk;
  assign mem_235_1_W0_data = W0_data[15:8];
  assign mem_235_1_W0_en = W0_en & W0_addr_sel == 8'heb;
  assign mem_235_1_W0_mask = W0_mask[1];
  assign mem_235_2_R0_addr = R0_addr[25:0];
  assign mem_235_2_R0_clk = R0_clk;
  assign mem_235_2_R0_en = R0_en & R0_addr_sel == 8'heb;
  assign mem_235_2_W0_addr = W0_addr[25:0];
  assign mem_235_2_W0_clk = W0_clk;
  assign mem_235_2_W0_data = W0_data[23:16];
  assign mem_235_2_W0_en = W0_en & W0_addr_sel == 8'heb;
  assign mem_235_2_W0_mask = W0_mask[2];
  assign mem_235_3_R0_addr = R0_addr[25:0];
  assign mem_235_3_R0_clk = R0_clk;
  assign mem_235_3_R0_en = R0_en & R0_addr_sel == 8'heb;
  assign mem_235_3_W0_addr = W0_addr[25:0];
  assign mem_235_3_W0_clk = W0_clk;
  assign mem_235_3_W0_data = W0_data[31:24];
  assign mem_235_3_W0_en = W0_en & W0_addr_sel == 8'heb;
  assign mem_235_3_W0_mask = W0_mask[3];
  assign mem_235_4_R0_addr = R0_addr[25:0];
  assign mem_235_4_R0_clk = R0_clk;
  assign mem_235_4_R0_en = R0_en & R0_addr_sel == 8'heb;
  assign mem_235_4_W0_addr = W0_addr[25:0];
  assign mem_235_4_W0_clk = W0_clk;
  assign mem_235_4_W0_data = W0_data[39:32];
  assign mem_235_4_W0_en = W0_en & W0_addr_sel == 8'heb;
  assign mem_235_4_W0_mask = W0_mask[4];
  assign mem_235_5_R0_addr = R0_addr[25:0];
  assign mem_235_5_R0_clk = R0_clk;
  assign mem_235_5_R0_en = R0_en & R0_addr_sel == 8'heb;
  assign mem_235_5_W0_addr = W0_addr[25:0];
  assign mem_235_5_W0_clk = W0_clk;
  assign mem_235_5_W0_data = W0_data[47:40];
  assign mem_235_5_W0_en = W0_en & W0_addr_sel == 8'heb;
  assign mem_235_5_W0_mask = W0_mask[5];
  assign mem_235_6_R0_addr = R0_addr[25:0];
  assign mem_235_6_R0_clk = R0_clk;
  assign mem_235_6_R0_en = R0_en & R0_addr_sel == 8'heb;
  assign mem_235_6_W0_addr = W0_addr[25:0];
  assign mem_235_6_W0_clk = W0_clk;
  assign mem_235_6_W0_data = W0_data[55:48];
  assign mem_235_6_W0_en = W0_en & W0_addr_sel == 8'heb;
  assign mem_235_6_W0_mask = W0_mask[6];
  assign mem_235_7_R0_addr = R0_addr[25:0];
  assign mem_235_7_R0_clk = R0_clk;
  assign mem_235_7_R0_en = R0_en & R0_addr_sel == 8'heb;
  assign mem_235_7_W0_addr = W0_addr[25:0];
  assign mem_235_7_W0_clk = W0_clk;
  assign mem_235_7_W0_data = W0_data[63:56];
  assign mem_235_7_W0_en = W0_en & W0_addr_sel == 8'heb;
  assign mem_235_7_W0_mask = W0_mask[7];
  assign mem_236_0_R0_addr = R0_addr[25:0];
  assign mem_236_0_R0_clk = R0_clk;
  assign mem_236_0_R0_en = R0_en & R0_addr_sel == 8'hec;
  assign mem_236_0_W0_addr = W0_addr[25:0];
  assign mem_236_0_W0_clk = W0_clk;
  assign mem_236_0_W0_data = W0_data[7:0];
  assign mem_236_0_W0_en = W0_en & W0_addr_sel == 8'hec;
  assign mem_236_0_W0_mask = W0_mask[0];
  assign mem_236_1_R0_addr = R0_addr[25:0];
  assign mem_236_1_R0_clk = R0_clk;
  assign mem_236_1_R0_en = R0_en & R0_addr_sel == 8'hec;
  assign mem_236_1_W0_addr = W0_addr[25:0];
  assign mem_236_1_W0_clk = W0_clk;
  assign mem_236_1_W0_data = W0_data[15:8];
  assign mem_236_1_W0_en = W0_en & W0_addr_sel == 8'hec;
  assign mem_236_1_W0_mask = W0_mask[1];
  assign mem_236_2_R0_addr = R0_addr[25:0];
  assign mem_236_2_R0_clk = R0_clk;
  assign mem_236_2_R0_en = R0_en & R0_addr_sel == 8'hec;
  assign mem_236_2_W0_addr = W0_addr[25:0];
  assign mem_236_2_W0_clk = W0_clk;
  assign mem_236_2_W0_data = W0_data[23:16];
  assign mem_236_2_W0_en = W0_en & W0_addr_sel == 8'hec;
  assign mem_236_2_W0_mask = W0_mask[2];
  assign mem_236_3_R0_addr = R0_addr[25:0];
  assign mem_236_3_R0_clk = R0_clk;
  assign mem_236_3_R0_en = R0_en & R0_addr_sel == 8'hec;
  assign mem_236_3_W0_addr = W0_addr[25:0];
  assign mem_236_3_W0_clk = W0_clk;
  assign mem_236_3_W0_data = W0_data[31:24];
  assign mem_236_3_W0_en = W0_en & W0_addr_sel == 8'hec;
  assign mem_236_3_W0_mask = W0_mask[3];
  assign mem_236_4_R0_addr = R0_addr[25:0];
  assign mem_236_4_R0_clk = R0_clk;
  assign mem_236_4_R0_en = R0_en & R0_addr_sel == 8'hec;
  assign mem_236_4_W0_addr = W0_addr[25:0];
  assign mem_236_4_W0_clk = W0_clk;
  assign mem_236_4_W0_data = W0_data[39:32];
  assign mem_236_4_W0_en = W0_en & W0_addr_sel == 8'hec;
  assign mem_236_4_W0_mask = W0_mask[4];
  assign mem_236_5_R0_addr = R0_addr[25:0];
  assign mem_236_5_R0_clk = R0_clk;
  assign mem_236_5_R0_en = R0_en & R0_addr_sel == 8'hec;
  assign mem_236_5_W0_addr = W0_addr[25:0];
  assign mem_236_5_W0_clk = W0_clk;
  assign mem_236_5_W0_data = W0_data[47:40];
  assign mem_236_5_W0_en = W0_en & W0_addr_sel == 8'hec;
  assign mem_236_5_W0_mask = W0_mask[5];
  assign mem_236_6_R0_addr = R0_addr[25:0];
  assign mem_236_6_R0_clk = R0_clk;
  assign mem_236_6_R0_en = R0_en & R0_addr_sel == 8'hec;
  assign mem_236_6_W0_addr = W0_addr[25:0];
  assign mem_236_6_W0_clk = W0_clk;
  assign mem_236_6_W0_data = W0_data[55:48];
  assign mem_236_6_W0_en = W0_en & W0_addr_sel == 8'hec;
  assign mem_236_6_W0_mask = W0_mask[6];
  assign mem_236_7_R0_addr = R0_addr[25:0];
  assign mem_236_7_R0_clk = R0_clk;
  assign mem_236_7_R0_en = R0_en & R0_addr_sel == 8'hec;
  assign mem_236_7_W0_addr = W0_addr[25:0];
  assign mem_236_7_W0_clk = W0_clk;
  assign mem_236_7_W0_data = W0_data[63:56];
  assign mem_236_7_W0_en = W0_en & W0_addr_sel == 8'hec;
  assign mem_236_7_W0_mask = W0_mask[7];
  assign mem_237_0_R0_addr = R0_addr[25:0];
  assign mem_237_0_R0_clk = R0_clk;
  assign mem_237_0_R0_en = R0_en & R0_addr_sel == 8'hed;
  assign mem_237_0_W0_addr = W0_addr[25:0];
  assign mem_237_0_W0_clk = W0_clk;
  assign mem_237_0_W0_data = W0_data[7:0];
  assign mem_237_0_W0_en = W0_en & W0_addr_sel == 8'hed;
  assign mem_237_0_W0_mask = W0_mask[0];
  assign mem_237_1_R0_addr = R0_addr[25:0];
  assign mem_237_1_R0_clk = R0_clk;
  assign mem_237_1_R0_en = R0_en & R0_addr_sel == 8'hed;
  assign mem_237_1_W0_addr = W0_addr[25:0];
  assign mem_237_1_W0_clk = W0_clk;
  assign mem_237_1_W0_data = W0_data[15:8];
  assign mem_237_1_W0_en = W0_en & W0_addr_sel == 8'hed;
  assign mem_237_1_W0_mask = W0_mask[1];
  assign mem_237_2_R0_addr = R0_addr[25:0];
  assign mem_237_2_R0_clk = R0_clk;
  assign mem_237_2_R0_en = R0_en & R0_addr_sel == 8'hed;
  assign mem_237_2_W0_addr = W0_addr[25:0];
  assign mem_237_2_W0_clk = W0_clk;
  assign mem_237_2_W0_data = W0_data[23:16];
  assign mem_237_2_W0_en = W0_en & W0_addr_sel == 8'hed;
  assign mem_237_2_W0_mask = W0_mask[2];
  assign mem_237_3_R0_addr = R0_addr[25:0];
  assign mem_237_3_R0_clk = R0_clk;
  assign mem_237_3_R0_en = R0_en & R0_addr_sel == 8'hed;
  assign mem_237_3_W0_addr = W0_addr[25:0];
  assign mem_237_3_W0_clk = W0_clk;
  assign mem_237_3_W0_data = W0_data[31:24];
  assign mem_237_3_W0_en = W0_en & W0_addr_sel == 8'hed;
  assign mem_237_3_W0_mask = W0_mask[3];
  assign mem_237_4_R0_addr = R0_addr[25:0];
  assign mem_237_4_R0_clk = R0_clk;
  assign mem_237_4_R0_en = R0_en & R0_addr_sel == 8'hed;
  assign mem_237_4_W0_addr = W0_addr[25:0];
  assign mem_237_4_W0_clk = W0_clk;
  assign mem_237_4_W0_data = W0_data[39:32];
  assign mem_237_4_W0_en = W0_en & W0_addr_sel == 8'hed;
  assign mem_237_4_W0_mask = W0_mask[4];
  assign mem_237_5_R0_addr = R0_addr[25:0];
  assign mem_237_5_R0_clk = R0_clk;
  assign mem_237_5_R0_en = R0_en & R0_addr_sel == 8'hed;
  assign mem_237_5_W0_addr = W0_addr[25:0];
  assign mem_237_5_W0_clk = W0_clk;
  assign mem_237_5_W0_data = W0_data[47:40];
  assign mem_237_5_W0_en = W0_en & W0_addr_sel == 8'hed;
  assign mem_237_5_W0_mask = W0_mask[5];
  assign mem_237_6_R0_addr = R0_addr[25:0];
  assign mem_237_6_R0_clk = R0_clk;
  assign mem_237_6_R0_en = R0_en & R0_addr_sel == 8'hed;
  assign mem_237_6_W0_addr = W0_addr[25:0];
  assign mem_237_6_W0_clk = W0_clk;
  assign mem_237_6_W0_data = W0_data[55:48];
  assign mem_237_6_W0_en = W0_en & W0_addr_sel == 8'hed;
  assign mem_237_6_W0_mask = W0_mask[6];
  assign mem_237_7_R0_addr = R0_addr[25:0];
  assign mem_237_7_R0_clk = R0_clk;
  assign mem_237_7_R0_en = R0_en & R0_addr_sel == 8'hed;
  assign mem_237_7_W0_addr = W0_addr[25:0];
  assign mem_237_7_W0_clk = W0_clk;
  assign mem_237_7_W0_data = W0_data[63:56];
  assign mem_237_7_W0_en = W0_en & W0_addr_sel == 8'hed;
  assign mem_237_7_W0_mask = W0_mask[7];
  assign mem_238_0_R0_addr = R0_addr[25:0];
  assign mem_238_0_R0_clk = R0_clk;
  assign mem_238_0_R0_en = R0_en & R0_addr_sel == 8'hee;
  assign mem_238_0_W0_addr = W0_addr[25:0];
  assign mem_238_0_W0_clk = W0_clk;
  assign mem_238_0_W0_data = W0_data[7:0];
  assign mem_238_0_W0_en = W0_en & W0_addr_sel == 8'hee;
  assign mem_238_0_W0_mask = W0_mask[0];
  assign mem_238_1_R0_addr = R0_addr[25:0];
  assign mem_238_1_R0_clk = R0_clk;
  assign mem_238_1_R0_en = R0_en & R0_addr_sel == 8'hee;
  assign mem_238_1_W0_addr = W0_addr[25:0];
  assign mem_238_1_W0_clk = W0_clk;
  assign mem_238_1_W0_data = W0_data[15:8];
  assign mem_238_1_W0_en = W0_en & W0_addr_sel == 8'hee;
  assign mem_238_1_W0_mask = W0_mask[1];
  assign mem_238_2_R0_addr = R0_addr[25:0];
  assign mem_238_2_R0_clk = R0_clk;
  assign mem_238_2_R0_en = R0_en & R0_addr_sel == 8'hee;
  assign mem_238_2_W0_addr = W0_addr[25:0];
  assign mem_238_2_W0_clk = W0_clk;
  assign mem_238_2_W0_data = W0_data[23:16];
  assign mem_238_2_W0_en = W0_en & W0_addr_sel == 8'hee;
  assign mem_238_2_W0_mask = W0_mask[2];
  assign mem_238_3_R0_addr = R0_addr[25:0];
  assign mem_238_3_R0_clk = R0_clk;
  assign mem_238_3_R0_en = R0_en & R0_addr_sel == 8'hee;
  assign mem_238_3_W0_addr = W0_addr[25:0];
  assign mem_238_3_W0_clk = W0_clk;
  assign mem_238_3_W0_data = W0_data[31:24];
  assign mem_238_3_W0_en = W0_en & W0_addr_sel == 8'hee;
  assign mem_238_3_W0_mask = W0_mask[3];
  assign mem_238_4_R0_addr = R0_addr[25:0];
  assign mem_238_4_R0_clk = R0_clk;
  assign mem_238_4_R0_en = R0_en & R0_addr_sel == 8'hee;
  assign mem_238_4_W0_addr = W0_addr[25:0];
  assign mem_238_4_W0_clk = W0_clk;
  assign mem_238_4_W0_data = W0_data[39:32];
  assign mem_238_4_W0_en = W0_en & W0_addr_sel == 8'hee;
  assign mem_238_4_W0_mask = W0_mask[4];
  assign mem_238_5_R0_addr = R0_addr[25:0];
  assign mem_238_5_R0_clk = R0_clk;
  assign mem_238_5_R0_en = R0_en & R0_addr_sel == 8'hee;
  assign mem_238_5_W0_addr = W0_addr[25:0];
  assign mem_238_5_W0_clk = W0_clk;
  assign mem_238_5_W0_data = W0_data[47:40];
  assign mem_238_5_W0_en = W0_en & W0_addr_sel == 8'hee;
  assign mem_238_5_W0_mask = W0_mask[5];
  assign mem_238_6_R0_addr = R0_addr[25:0];
  assign mem_238_6_R0_clk = R0_clk;
  assign mem_238_6_R0_en = R0_en & R0_addr_sel == 8'hee;
  assign mem_238_6_W0_addr = W0_addr[25:0];
  assign mem_238_6_W0_clk = W0_clk;
  assign mem_238_6_W0_data = W0_data[55:48];
  assign mem_238_6_W0_en = W0_en & W0_addr_sel == 8'hee;
  assign mem_238_6_W0_mask = W0_mask[6];
  assign mem_238_7_R0_addr = R0_addr[25:0];
  assign mem_238_7_R0_clk = R0_clk;
  assign mem_238_7_R0_en = R0_en & R0_addr_sel == 8'hee;
  assign mem_238_7_W0_addr = W0_addr[25:0];
  assign mem_238_7_W0_clk = W0_clk;
  assign mem_238_7_W0_data = W0_data[63:56];
  assign mem_238_7_W0_en = W0_en & W0_addr_sel == 8'hee;
  assign mem_238_7_W0_mask = W0_mask[7];
  assign mem_239_0_R0_addr = R0_addr[25:0];
  assign mem_239_0_R0_clk = R0_clk;
  assign mem_239_0_R0_en = R0_en & R0_addr_sel == 8'hef;
  assign mem_239_0_W0_addr = W0_addr[25:0];
  assign mem_239_0_W0_clk = W0_clk;
  assign mem_239_0_W0_data = W0_data[7:0];
  assign mem_239_0_W0_en = W0_en & W0_addr_sel == 8'hef;
  assign mem_239_0_W0_mask = W0_mask[0];
  assign mem_239_1_R0_addr = R0_addr[25:0];
  assign mem_239_1_R0_clk = R0_clk;
  assign mem_239_1_R0_en = R0_en & R0_addr_sel == 8'hef;
  assign mem_239_1_W0_addr = W0_addr[25:0];
  assign mem_239_1_W0_clk = W0_clk;
  assign mem_239_1_W0_data = W0_data[15:8];
  assign mem_239_1_W0_en = W0_en & W0_addr_sel == 8'hef;
  assign mem_239_1_W0_mask = W0_mask[1];
  assign mem_239_2_R0_addr = R0_addr[25:0];
  assign mem_239_2_R0_clk = R0_clk;
  assign mem_239_2_R0_en = R0_en & R0_addr_sel == 8'hef;
  assign mem_239_2_W0_addr = W0_addr[25:0];
  assign mem_239_2_W0_clk = W0_clk;
  assign mem_239_2_W0_data = W0_data[23:16];
  assign mem_239_2_W0_en = W0_en & W0_addr_sel == 8'hef;
  assign mem_239_2_W0_mask = W0_mask[2];
  assign mem_239_3_R0_addr = R0_addr[25:0];
  assign mem_239_3_R0_clk = R0_clk;
  assign mem_239_3_R0_en = R0_en & R0_addr_sel == 8'hef;
  assign mem_239_3_W0_addr = W0_addr[25:0];
  assign mem_239_3_W0_clk = W0_clk;
  assign mem_239_3_W0_data = W0_data[31:24];
  assign mem_239_3_W0_en = W0_en & W0_addr_sel == 8'hef;
  assign mem_239_3_W0_mask = W0_mask[3];
  assign mem_239_4_R0_addr = R0_addr[25:0];
  assign mem_239_4_R0_clk = R0_clk;
  assign mem_239_4_R0_en = R0_en & R0_addr_sel == 8'hef;
  assign mem_239_4_W0_addr = W0_addr[25:0];
  assign mem_239_4_W0_clk = W0_clk;
  assign mem_239_4_W0_data = W0_data[39:32];
  assign mem_239_4_W0_en = W0_en & W0_addr_sel == 8'hef;
  assign mem_239_4_W0_mask = W0_mask[4];
  assign mem_239_5_R0_addr = R0_addr[25:0];
  assign mem_239_5_R0_clk = R0_clk;
  assign mem_239_5_R0_en = R0_en & R0_addr_sel == 8'hef;
  assign mem_239_5_W0_addr = W0_addr[25:0];
  assign mem_239_5_W0_clk = W0_clk;
  assign mem_239_5_W0_data = W0_data[47:40];
  assign mem_239_5_W0_en = W0_en & W0_addr_sel == 8'hef;
  assign mem_239_5_W0_mask = W0_mask[5];
  assign mem_239_6_R0_addr = R0_addr[25:0];
  assign mem_239_6_R0_clk = R0_clk;
  assign mem_239_6_R0_en = R0_en & R0_addr_sel == 8'hef;
  assign mem_239_6_W0_addr = W0_addr[25:0];
  assign mem_239_6_W0_clk = W0_clk;
  assign mem_239_6_W0_data = W0_data[55:48];
  assign mem_239_6_W0_en = W0_en & W0_addr_sel == 8'hef;
  assign mem_239_6_W0_mask = W0_mask[6];
  assign mem_239_7_R0_addr = R0_addr[25:0];
  assign mem_239_7_R0_clk = R0_clk;
  assign mem_239_7_R0_en = R0_en & R0_addr_sel == 8'hef;
  assign mem_239_7_W0_addr = W0_addr[25:0];
  assign mem_239_7_W0_clk = W0_clk;
  assign mem_239_7_W0_data = W0_data[63:56];
  assign mem_239_7_W0_en = W0_en & W0_addr_sel == 8'hef;
  assign mem_239_7_W0_mask = W0_mask[7];
  assign mem_240_0_R0_addr = R0_addr[25:0];
  assign mem_240_0_R0_clk = R0_clk;
  assign mem_240_0_R0_en = R0_en & R0_addr_sel == 8'hf0;
  assign mem_240_0_W0_addr = W0_addr[25:0];
  assign mem_240_0_W0_clk = W0_clk;
  assign mem_240_0_W0_data = W0_data[7:0];
  assign mem_240_0_W0_en = W0_en & W0_addr_sel == 8'hf0;
  assign mem_240_0_W0_mask = W0_mask[0];
  assign mem_240_1_R0_addr = R0_addr[25:0];
  assign mem_240_1_R0_clk = R0_clk;
  assign mem_240_1_R0_en = R0_en & R0_addr_sel == 8'hf0;
  assign mem_240_1_W0_addr = W0_addr[25:0];
  assign mem_240_1_W0_clk = W0_clk;
  assign mem_240_1_W0_data = W0_data[15:8];
  assign mem_240_1_W0_en = W0_en & W0_addr_sel == 8'hf0;
  assign mem_240_1_W0_mask = W0_mask[1];
  assign mem_240_2_R0_addr = R0_addr[25:0];
  assign mem_240_2_R0_clk = R0_clk;
  assign mem_240_2_R0_en = R0_en & R0_addr_sel == 8'hf0;
  assign mem_240_2_W0_addr = W0_addr[25:0];
  assign mem_240_2_W0_clk = W0_clk;
  assign mem_240_2_W0_data = W0_data[23:16];
  assign mem_240_2_W0_en = W0_en & W0_addr_sel == 8'hf0;
  assign mem_240_2_W0_mask = W0_mask[2];
  assign mem_240_3_R0_addr = R0_addr[25:0];
  assign mem_240_3_R0_clk = R0_clk;
  assign mem_240_3_R0_en = R0_en & R0_addr_sel == 8'hf0;
  assign mem_240_3_W0_addr = W0_addr[25:0];
  assign mem_240_3_W0_clk = W0_clk;
  assign mem_240_3_W0_data = W0_data[31:24];
  assign mem_240_3_W0_en = W0_en & W0_addr_sel == 8'hf0;
  assign mem_240_3_W0_mask = W0_mask[3];
  assign mem_240_4_R0_addr = R0_addr[25:0];
  assign mem_240_4_R0_clk = R0_clk;
  assign mem_240_4_R0_en = R0_en & R0_addr_sel == 8'hf0;
  assign mem_240_4_W0_addr = W0_addr[25:0];
  assign mem_240_4_W0_clk = W0_clk;
  assign mem_240_4_W0_data = W0_data[39:32];
  assign mem_240_4_W0_en = W0_en & W0_addr_sel == 8'hf0;
  assign mem_240_4_W0_mask = W0_mask[4];
  assign mem_240_5_R0_addr = R0_addr[25:0];
  assign mem_240_5_R0_clk = R0_clk;
  assign mem_240_5_R0_en = R0_en & R0_addr_sel == 8'hf0;
  assign mem_240_5_W0_addr = W0_addr[25:0];
  assign mem_240_5_W0_clk = W0_clk;
  assign mem_240_5_W0_data = W0_data[47:40];
  assign mem_240_5_W0_en = W0_en & W0_addr_sel == 8'hf0;
  assign mem_240_5_W0_mask = W0_mask[5];
  assign mem_240_6_R0_addr = R0_addr[25:0];
  assign mem_240_6_R0_clk = R0_clk;
  assign mem_240_6_R0_en = R0_en & R0_addr_sel == 8'hf0;
  assign mem_240_6_W0_addr = W0_addr[25:0];
  assign mem_240_6_W0_clk = W0_clk;
  assign mem_240_6_W0_data = W0_data[55:48];
  assign mem_240_6_W0_en = W0_en & W0_addr_sel == 8'hf0;
  assign mem_240_6_W0_mask = W0_mask[6];
  assign mem_240_7_R0_addr = R0_addr[25:0];
  assign mem_240_7_R0_clk = R0_clk;
  assign mem_240_7_R0_en = R0_en & R0_addr_sel == 8'hf0;
  assign mem_240_7_W0_addr = W0_addr[25:0];
  assign mem_240_7_W0_clk = W0_clk;
  assign mem_240_7_W0_data = W0_data[63:56];
  assign mem_240_7_W0_en = W0_en & W0_addr_sel == 8'hf0;
  assign mem_240_7_W0_mask = W0_mask[7];
  assign mem_241_0_R0_addr = R0_addr[25:0];
  assign mem_241_0_R0_clk = R0_clk;
  assign mem_241_0_R0_en = R0_en & R0_addr_sel == 8'hf1;
  assign mem_241_0_W0_addr = W0_addr[25:0];
  assign mem_241_0_W0_clk = W0_clk;
  assign mem_241_0_W0_data = W0_data[7:0];
  assign mem_241_0_W0_en = W0_en & W0_addr_sel == 8'hf1;
  assign mem_241_0_W0_mask = W0_mask[0];
  assign mem_241_1_R0_addr = R0_addr[25:0];
  assign mem_241_1_R0_clk = R0_clk;
  assign mem_241_1_R0_en = R0_en & R0_addr_sel == 8'hf1;
  assign mem_241_1_W0_addr = W0_addr[25:0];
  assign mem_241_1_W0_clk = W0_clk;
  assign mem_241_1_W0_data = W0_data[15:8];
  assign mem_241_1_W0_en = W0_en & W0_addr_sel == 8'hf1;
  assign mem_241_1_W0_mask = W0_mask[1];
  assign mem_241_2_R0_addr = R0_addr[25:0];
  assign mem_241_2_R0_clk = R0_clk;
  assign mem_241_2_R0_en = R0_en & R0_addr_sel == 8'hf1;
  assign mem_241_2_W0_addr = W0_addr[25:0];
  assign mem_241_2_W0_clk = W0_clk;
  assign mem_241_2_W0_data = W0_data[23:16];
  assign mem_241_2_W0_en = W0_en & W0_addr_sel == 8'hf1;
  assign mem_241_2_W0_mask = W0_mask[2];
  assign mem_241_3_R0_addr = R0_addr[25:0];
  assign mem_241_3_R0_clk = R0_clk;
  assign mem_241_3_R0_en = R0_en & R0_addr_sel == 8'hf1;
  assign mem_241_3_W0_addr = W0_addr[25:0];
  assign mem_241_3_W0_clk = W0_clk;
  assign mem_241_3_W0_data = W0_data[31:24];
  assign mem_241_3_W0_en = W0_en & W0_addr_sel == 8'hf1;
  assign mem_241_3_W0_mask = W0_mask[3];
  assign mem_241_4_R0_addr = R0_addr[25:0];
  assign mem_241_4_R0_clk = R0_clk;
  assign mem_241_4_R0_en = R0_en & R0_addr_sel == 8'hf1;
  assign mem_241_4_W0_addr = W0_addr[25:0];
  assign mem_241_4_W0_clk = W0_clk;
  assign mem_241_4_W0_data = W0_data[39:32];
  assign mem_241_4_W0_en = W0_en & W0_addr_sel == 8'hf1;
  assign mem_241_4_W0_mask = W0_mask[4];
  assign mem_241_5_R0_addr = R0_addr[25:0];
  assign mem_241_5_R0_clk = R0_clk;
  assign mem_241_5_R0_en = R0_en & R0_addr_sel == 8'hf1;
  assign mem_241_5_W0_addr = W0_addr[25:0];
  assign mem_241_5_W0_clk = W0_clk;
  assign mem_241_5_W0_data = W0_data[47:40];
  assign mem_241_5_W0_en = W0_en & W0_addr_sel == 8'hf1;
  assign mem_241_5_W0_mask = W0_mask[5];
  assign mem_241_6_R0_addr = R0_addr[25:0];
  assign mem_241_6_R0_clk = R0_clk;
  assign mem_241_6_R0_en = R0_en & R0_addr_sel == 8'hf1;
  assign mem_241_6_W0_addr = W0_addr[25:0];
  assign mem_241_6_W0_clk = W0_clk;
  assign mem_241_6_W0_data = W0_data[55:48];
  assign mem_241_6_W0_en = W0_en & W0_addr_sel == 8'hf1;
  assign mem_241_6_W0_mask = W0_mask[6];
  assign mem_241_7_R0_addr = R0_addr[25:0];
  assign mem_241_7_R0_clk = R0_clk;
  assign mem_241_7_R0_en = R0_en & R0_addr_sel == 8'hf1;
  assign mem_241_7_W0_addr = W0_addr[25:0];
  assign mem_241_7_W0_clk = W0_clk;
  assign mem_241_7_W0_data = W0_data[63:56];
  assign mem_241_7_W0_en = W0_en & W0_addr_sel == 8'hf1;
  assign mem_241_7_W0_mask = W0_mask[7];
  assign mem_242_0_R0_addr = R0_addr[25:0];
  assign mem_242_0_R0_clk = R0_clk;
  assign mem_242_0_R0_en = R0_en & R0_addr_sel == 8'hf2;
  assign mem_242_0_W0_addr = W0_addr[25:0];
  assign mem_242_0_W0_clk = W0_clk;
  assign mem_242_0_W0_data = W0_data[7:0];
  assign mem_242_0_W0_en = W0_en & W0_addr_sel == 8'hf2;
  assign mem_242_0_W0_mask = W0_mask[0];
  assign mem_242_1_R0_addr = R0_addr[25:0];
  assign mem_242_1_R0_clk = R0_clk;
  assign mem_242_1_R0_en = R0_en & R0_addr_sel == 8'hf2;
  assign mem_242_1_W0_addr = W0_addr[25:0];
  assign mem_242_1_W0_clk = W0_clk;
  assign mem_242_1_W0_data = W0_data[15:8];
  assign mem_242_1_W0_en = W0_en & W0_addr_sel == 8'hf2;
  assign mem_242_1_W0_mask = W0_mask[1];
  assign mem_242_2_R0_addr = R0_addr[25:0];
  assign mem_242_2_R0_clk = R0_clk;
  assign mem_242_2_R0_en = R0_en & R0_addr_sel == 8'hf2;
  assign mem_242_2_W0_addr = W0_addr[25:0];
  assign mem_242_2_W0_clk = W0_clk;
  assign mem_242_2_W0_data = W0_data[23:16];
  assign mem_242_2_W0_en = W0_en & W0_addr_sel == 8'hf2;
  assign mem_242_2_W0_mask = W0_mask[2];
  assign mem_242_3_R0_addr = R0_addr[25:0];
  assign mem_242_3_R0_clk = R0_clk;
  assign mem_242_3_R0_en = R0_en & R0_addr_sel == 8'hf2;
  assign mem_242_3_W0_addr = W0_addr[25:0];
  assign mem_242_3_W0_clk = W0_clk;
  assign mem_242_3_W0_data = W0_data[31:24];
  assign mem_242_3_W0_en = W0_en & W0_addr_sel == 8'hf2;
  assign mem_242_3_W0_mask = W0_mask[3];
  assign mem_242_4_R0_addr = R0_addr[25:0];
  assign mem_242_4_R0_clk = R0_clk;
  assign mem_242_4_R0_en = R0_en & R0_addr_sel == 8'hf2;
  assign mem_242_4_W0_addr = W0_addr[25:0];
  assign mem_242_4_W0_clk = W0_clk;
  assign mem_242_4_W0_data = W0_data[39:32];
  assign mem_242_4_W0_en = W0_en & W0_addr_sel == 8'hf2;
  assign mem_242_4_W0_mask = W0_mask[4];
  assign mem_242_5_R0_addr = R0_addr[25:0];
  assign mem_242_5_R0_clk = R0_clk;
  assign mem_242_5_R0_en = R0_en & R0_addr_sel == 8'hf2;
  assign mem_242_5_W0_addr = W0_addr[25:0];
  assign mem_242_5_W0_clk = W0_clk;
  assign mem_242_5_W0_data = W0_data[47:40];
  assign mem_242_5_W0_en = W0_en & W0_addr_sel == 8'hf2;
  assign mem_242_5_W0_mask = W0_mask[5];
  assign mem_242_6_R0_addr = R0_addr[25:0];
  assign mem_242_6_R0_clk = R0_clk;
  assign mem_242_6_R0_en = R0_en & R0_addr_sel == 8'hf2;
  assign mem_242_6_W0_addr = W0_addr[25:0];
  assign mem_242_6_W0_clk = W0_clk;
  assign mem_242_6_W0_data = W0_data[55:48];
  assign mem_242_6_W0_en = W0_en & W0_addr_sel == 8'hf2;
  assign mem_242_6_W0_mask = W0_mask[6];
  assign mem_242_7_R0_addr = R0_addr[25:0];
  assign mem_242_7_R0_clk = R0_clk;
  assign mem_242_7_R0_en = R0_en & R0_addr_sel == 8'hf2;
  assign mem_242_7_W0_addr = W0_addr[25:0];
  assign mem_242_7_W0_clk = W0_clk;
  assign mem_242_7_W0_data = W0_data[63:56];
  assign mem_242_7_W0_en = W0_en & W0_addr_sel == 8'hf2;
  assign mem_242_7_W0_mask = W0_mask[7];
  assign mem_243_0_R0_addr = R0_addr[25:0];
  assign mem_243_0_R0_clk = R0_clk;
  assign mem_243_0_R0_en = R0_en & R0_addr_sel == 8'hf3;
  assign mem_243_0_W0_addr = W0_addr[25:0];
  assign mem_243_0_W0_clk = W0_clk;
  assign mem_243_0_W0_data = W0_data[7:0];
  assign mem_243_0_W0_en = W0_en & W0_addr_sel == 8'hf3;
  assign mem_243_0_W0_mask = W0_mask[0];
  assign mem_243_1_R0_addr = R0_addr[25:0];
  assign mem_243_1_R0_clk = R0_clk;
  assign mem_243_1_R0_en = R0_en & R0_addr_sel == 8'hf3;
  assign mem_243_1_W0_addr = W0_addr[25:0];
  assign mem_243_1_W0_clk = W0_clk;
  assign mem_243_1_W0_data = W0_data[15:8];
  assign mem_243_1_W0_en = W0_en & W0_addr_sel == 8'hf3;
  assign mem_243_1_W0_mask = W0_mask[1];
  assign mem_243_2_R0_addr = R0_addr[25:0];
  assign mem_243_2_R0_clk = R0_clk;
  assign mem_243_2_R0_en = R0_en & R0_addr_sel == 8'hf3;
  assign mem_243_2_W0_addr = W0_addr[25:0];
  assign mem_243_2_W0_clk = W0_clk;
  assign mem_243_2_W0_data = W0_data[23:16];
  assign mem_243_2_W0_en = W0_en & W0_addr_sel == 8'hf3;
  assign mem_243_2_W0_mask = W0_mask[2];
  assign mem_243_3_R0_addr = R0_addr[25:0];
  assign mem_243_3_R0_clk = R0_clk;
  assign mem_243_3_R0_en = R0_en & R0_addr_sel == 8'hf3;
  assign mem_243_3_W0_addr = W0_addr[25:0];
  assign mem_243_3_W0_clk = W0_clk;
  assign mem_243_3_W0_data = W0_data[31:24];
  assign mem_243_3_W0_en = W0_en & W0_addr_sel == 8'hf3;
  assign mem_243_3_W0_mask = W0_mask[3];
  assign mem_243_4_R0_addr = R0_addr[25:0];
  assign mem_243_4_R0_clk = R0_clk;
  assign mem_243_4_R0_en = R0_en & R0_addr_sel == 8'hf3;
  assign mem_243_4_W0_addr = W0_addr[25:0];
  assign mem_243_4_W0_clk = W0_clk;
  assign mem_243_4_W0_data = W0_data[39:32];
  assign mem_243_4_W0_en = W0_en & W0_addr_sel == 8'hf3;
  assign mem_243_4_W0_mask = W0_mask[4];
  assign mem_243_5_R0_addr = R0_addr[25:0];
  assign mem_243_5_R0_clk = R0_clk;
  assign mem_243_5_R0_en = R0_en & R0_addr_sel == 8'hf3;
  assign mem_243_5_W0_addr = W0_addr[25:0];
  assign mem_243_5_W0_clk = W0_clk;
  assign mem_243_5_W0_data = W0_data[47:40];
  assign mem_243_5_W0_en = W0_en & W0_addr_sel == 8'hf3;
  assign mem_243_5_W0_mask = W0_mask[5];
  assign mem_243_6_R0_addr = R0_addr[25:0];
  assign mem_243_6_R0_clk = R0_clk;
  assign mem_243_6_R0_en = R0_en & R0_addr_sel == 8'hf3;
  assign mem_243_6_W0_addr = W0_addr[25:0];
  assign mem_243_6_W0_clk = W0_clk;
  assign mem_243_6_W0_data = W0_data[55:48];
  assign mem_243_6_W0_en = W0_en & W0_addr_sel == 8'hf3;
  assign mem_243_6_W0_mask = W0_mask[6];
  assign mem_243_7_R0_addr = R0_addr[25:0];
  assign mem_243_7_R0_clk = R0_clk;
  assign mem_243_7_R0_en = R0_en & R0_addr_sel == 8'hf3;
  assign mem_243_7_W0_addr = W0_addr[25:0];
  assign mem_243_7_W0_clk = W0_clk;
  assign mem_243_7_W0_data = W0_data[63:56];
  assign mem_243_7_W0_en = W0_en & W0_addr_sel == 8'hf3;
  assign mem_243_7_W0_mask = W0_mask[7];
  assign mem_244_0_R0_addr = R0_addr[25:0];
  assign mem_244_0_R0_clk = R0_clk;
  assign mem_244_0_R0_en = R0_en & R0_addr_sel == 8'hf4;
  assign mem_244_0_W0_addr = W0_addr[25:0];
  assign mem_244_0_W0_clk = W0_clk;
  assign mem_244_0_W0_data = W0_data[7:0];
  assign mem_244_0_W0_en = W0_en & W0_addr_sel == 8'hf4;
  assign mem_244_0_W0_mask = W0_mask[0];
  assign mem_244_1_R0_addr = R0_addr[25:0];
  assign mem_244_1_R0_clk = R0_clk;
  assign mem_244_1_R0_en = R0_en & R0_addr_sel == 8'hf4;
  assign mem_244_1_W0_addr = W0_addr[25:0];
  assign mem_244_1_W0_clk = W0_clk;
  assign mem_244_1_W0_data = W0_data[15:8];
  assign mem_244_1_W0_en = W0_en & W0_addr_sel == 8'hf4;
  assign mem_244_1_W0_mask = W0_mask[1];
  assign mem_244_2_R0_addr = R0_addr[25:0];
  assign mem_244_2_R0_clk = R0_clk;
  assign mem_244_2_R0_en = R0_en & R0_addr_sel == 8'hf4;
  assign mem_244_2_W0_addr = W0_addr[25:0];
  assign mem_244_2_W0_clk = W0_clk;
  assign mem_244_2_W0_data = W0_data[23:16];
  assign mem_244_2_W0_en = W0_en & W0_addr_sel == 8'hf4;
  assign mem_244_2_W0_mask = W0_mask[2];
  assign mem_244_3_R0_addr = R0_addr[25:0];
  assign mem_244_3_R0_clk = R0_clk;
  assign mem_244_3_R0_en = R0_en & R0_addr_sel == 8'hf4;
  assign mem_244_3_W0_addr = W0_addr[25:0];
  assign mem_244_3_W0_clk = W0_clk;
  assign mem_244_3_W0_data = W0_data[31:24];
  assign mem_244_3_W0_en = W0_en & W0_addr_sel == 8'hf4;
  assign mem_244_3_W0_mask = W0_mask[3];
  assign mem_244_4_R0_addr = R0_addr[25:0];
  assign mem_244_4_R0_clk = R0_clk;
  assign mem_244_4_R0_en = R0_en & R0_addr_sel == 8'hf4;
  assign mem_244_4_W0_addr = W0_addr[25:0];
  assign mem_244_4_W0_clk = W0_clk;
  assign mem_244_4_W0_data = W0_data[39:32];
  assign mem_244_4_W0_en = W0_en & W0_addr_sel == 8'hf4;
  assign mem_244_4_W0_mask = W0_mask[4];
  assign mem_244_5_R0_addr = R0_addr[25:0];
  assign mem_244_5_R0_clk = R0_clk;
  assign mem_244_5_R0_en = R0_en & R0_addr_sel == 8'hf4;
  assign mem_244_5_W0_addr = W0_addr[25:0];
  assign mem_244_5_W0_clk = W0_clk;
  assign mem_244_5_W0_data = W0_data[47:40];
  assign mem_244_5_W0_en = W0_en & W0_addr_sel == 8'hf4;
  assign mem_244_5_W0_mask = W0_mask[5];
  assign mem_244_6_R0_addr = R0_addr[25:0];
  assign mem_244_6_R0_clk = R0_clk;
  assign mem_244_6_R0_en = R0_en & R0_addr_sel == 8'hf4;
  assign mem_244_6_W0_addr = W0_addr[25:0];
  assign mem_244_6_W0_clk = W0_clk;
  assign mem_244_6_W0_data = W0_data[55:48];
  assign mem_244_6_W0_en = W0_en & W0_addr_sel == 8'hf4;
  assign mem_244_6_W0_mask = W0_mask[6];
  assign mem_244_7_R0_addr = R0_addr[25:0];
  assign mem_244_7_R0_clk = R0_clk;
  assign mem_244_7_R0_en = R0_en & R0_addr_sel == 8'hf4;
  assign mem_244_7_W0_addr = W0_addr[25:0];
  assign mem_244_7_W0_clk = W0_clk;
  assign mem_244_7_W0_data = W0_data[63:56];
  assign mem_244_7_W0_en = W0_en & W0_addr_sel == 8'hf4;
  assign mem_244_7_W0_mask = W0_mask[7];
  assign mem_245_0_R0_addr = R0_addr[25:0];
  assign mem_245_0_R0_clk = R0_clk;
  assign mem_245_0_R0_en = R0_en & R0_addr_sel == 8'hf5;
  assign mem_245_0_W0_addr = W0_addr[25:0];
  assign mem_245_0_W0_clk = W0_clk;
  assign mem_245_0_W0_data = W0_data[7:0];
  assign mem_245_0_W0_en = W0_en & W0_addr_sel == 8'hf5;
  assign mem_245_0_W0_mask = W0_mask[0];
  assign mem_245_1_R0_addr = R0_addr[25:0];
  assign mem_245_1_R0_clk = R0_clk;
  assign mem_245_1_R0_en = R0_en & R0_addr_sel == 8'hf5;
  assign mem_245_1_W0_addr = W0_addr[25:0];
  assign mem_245_1_W0_clk = W0_clk;
  assign mem_245_1_W0_data = W0_data[15:8];
  assign mem_245_1_W0_en = W0_en & W0_addr_sel == 8'hf5;
  assign mem_245_1_W0_mask = W0_mask[1];
  assign mem_245_2_R0_addr = R0_addr[25:0];
  assign mem_245_2_R0_clk = R0_clk;
  assign mem_245_2_R0_en = R0_en & R0_addr_sel == 8'hf5;
  assign mem_245_2_W0_addr = W0_addr[25:0];
  assign mem_245_2_W0_clk = W0_clk;
  assign mem_245_2_W0_data = W0_data[23:16];
  assign mem_245_2_W0_en = W0_en & W0_addr_sel == 8'hf5;
  assign mem_245_2_W0_mask = W0_mask[2];
  assign mem_245_3_R0_addr = R0_addr[25:0];
  assign mem_245_3_R0_clk = R0_clk;
  assign mem_245_3_R0_en = R0_en & R0_addr_sel == 8'hf5;
  assign mem_245_3_W0_addr = W0_addr[25:0];
  assign mem_245_3_W0_clk = W0_clk;
  assign mem_245_3_W0_data = W0_data[31:24];
  assign mem_245_3_W0_en = W0_en & W0_addr_sel == 8'hf5;
  assign mem_245_3_W0_mask = W0_mask[3];
  assign mem_245_4_R0_addr = R0_addr[25:0];
  assign mem_245_4_R0_clk = R0_clk;
  assign mem_245_4_R0_en = R0_en & R0_addr_sel == 8'hf5;
  assign mem_245_4_W0_addr = W0_addr[25:0];
  assign mem_245_4_W0_clk = W0_clk;
  assign mem_245_4_W0_data = W0_data[39:32];
  assign mem_245_4_W0_en = W0_en & W0_addr_sel == 8'hf5;
  assign mem_245_4_W0_mask = W0_mask[4];
  assign mem_245_5_R0_addr = R0_addr[25:0];
  assign mem_245_5_R0_clk = R0_clk;
  assign mem_245_5_R0_en = R0_en & R0_addr_sel == 8'hf5;
  assign mem_245_5_W0_addr = W0_addr[25:0];
  assign mem_245_5_W0_clk = W0_clk;
  assign mem_245_5_W0_data = W0_data[47:40];
  assign mem_245_5_W0_en = W0_en & W0_addr_sel == 8'hf5;
  assign mem_245_5_W0_mask = W0_mask[5];
  assign mem_245_6_R0_addr = R0_addr[25:0];
  assign mem_245_6_R0_clk = R0_clk;
  assign mem_245_6_R0_en = R0_en & R0_addr_sel == 8'hf5;
  assign mem_245_6_W0_addr = W0_addr[25:0];
  assign mem_245_6_W0_clk = W0_clk;
  assign mem_245_6_W0_data = W0_data[55:48];
  assign mem_245_6_W0_en = W0_en & W0_addr_sel == 8'hf5;
  assign mem_245_6_W0_mask = W0_mask[6];
  assign mem_245_7_R0_addr = R0_addr[25:0];
  assign mem_245_7_R0_clk = R0_clk;
  assign mem_245_7_R0_en = R0_en & R0_addr_sel == 8'hf5;
  assign mem_245_7_W0_addr = W0_addr[25:0];
  assign mem_245_7_W0_clk = W0_clk;
  assign mem_245_7_W0_data = W0_data[63:56];
  assign mem_245_7_W0_en = W0_en & W0_addr_sel == 8'hf5;
  assign mem_245_7_W0_mask = W0_mask[7];
  assign mem_246_0_R0_addr = R0_addr[25:0];
  assign mem_246_0_R0_clk = R0_clk;
  assign mem_246_0_R0_en = R0_en & R0_addr_sel == 8'hf6;
  assign mem_246_0_W0_addr = W0_addr[25:0];
  assign mem_246_0_W0_clk = W0_clk;
  assign mem_246_0_W0_data = W0_data[7:0];
  assign mem_246_0_W0_en = W0_en & W0_addr_sel == 8'hf6;
  assign mem_246_0_W0_mask = W0_mask[0];
  assign mem_246_1_R0_addr = R0_addr[25:0];
  assign mem_246_1_R0_clk = R0_clk;
  assign mem_246_1_R0_en = R0_en & R0_addr_sel == 8'hf6;
  assign mem_246_1_W0_addr = W0_addr[25:0];
  assign mem_246_1_W0_clk = W0_clk;
  assign mem_246_1_W0_data = W0_data[15:8];
  assign mem_246_1_W0_en = W0_en & W0_addr_sel == 8'hf6;
  assign mem_246_1_W0_mask = W0_mask[1];
  assign mem_246_2_R0_addr = R0_addr[25:0];
  assign mem_246_2_R0_clk = R0_clk;
  assign mem_246_2_R0_en = R0_en & R0_addr_sel == 8'hf6;
  assign mem_246_2_W0_addr = W0_addr[25:0];
  assign mem_246_2_W0_clk = W0_clk;
  assign mem_246_2_W0_data = W0_data[23:16];
  assign mem_246_2_W0_en = W0_en & W0_addr_sel == 8'hf6;
  assign mem_246_2_W0_mask = W0_mask[2];
  assign mem_246_3_R0_addr = R0_addr[25:0];
  assign mem_246_3_R0_clk = R0_clk;
  assign mem_246_3_R0_en = R0_en & R0_addr_sel == 8'hf6;
  assign mem_246_3_W0_addr = W0_addr[25:0];
  assign mem_246_3_W0_clk = W0_clk;
  assign mem_246_3_W0_data = W0_data[31:24];
  assign mem_246_3_W0_en = W0_en & W0_addr_sel == 8'hf6;
  assign mem_246_3_W0_mask = W0_mask[3];
  assign mem_246_4_R0_addr = R0_addr[25:0];
  assign mem_246_4_R0_clk = R0_clk;
  assign mem_246_4_R0_en = R0_en & R0_addr_sel == 8'hf6;
  assign mem_246_4_W0_addr = W0_addr[25:0];
  assign mem_246_4_W0_clk = W0_clk;
  assign mem_246_4_W0_data = W0_data[39:32];
  assign mem_246_4_W0_en = W0_en & W0_addr_sel == 8'hf6;
  assign mem_246_4_W0_mask = W0_mask[4];
  assign mem_246_5_R0_addr = R0_addr[25:0];
  assign mem_246_5_R0_clk = R0_clk;
  assign mem_246_5_R0_en = R0_en & R0_addr_sel == 8'hf6;
  assign mem_246_5_W0_addr = W0_addr[25:0];
  assign mem_246_5_W0_clk = W0_clk;
  assign mem_246_5_W0_data = W0_data[47:40];
  assign mem_246_5_W0_en = W0_en & W0_addr_sel == 8'hf6;
  assign mem_246_5_W0_mask = W0_mask[5];
  assign mem_246_6_R0_addr = R0_addr[25:0];
  assign mem_246_6_R0_clk = R0_clk;
  assign mem_246_6_R0_en = R0_en & R0_addr_sel == 8'hf6;
  assign mem_246_6_W0_addr = W0_addr[25:0];
  assign mem_246_6_W0_clk = W0_clk;
  assign mem_246_6_W0_data = W0_data[55:48];
  assign mem_246_6_W0_en = W0_en & W0_addr_sel == 8'hf6;
  assign mem_246_6_W0_mask = W0_mask[6];
  assign mem_246_7_R0_addr = R0_addr[25:0];
  assign mem_246_7_R0_clk = R0_clk;
  assign mem_246_7_R0_en = R0_en & R0_addr_sel == 8'hf6;
  assign mem_246_7_W0_addr = W0_addr[25:0];
  assign mem_246_7_W0_clk = W0_clk;
  assign mem_246_7_W0_data = W0_data[63:56];
  assign mem_246_7_W0_en = W0_en & W0_addr_sel == 8'hf6;
  assign mem_246_7_W0_mask = W0_mask[7];
  assign mem_247_0_R0_addr = R0_addr[25:0];
  assign mem_247_0_R0_clk = R0_clk;
  assign mem_247_0_R0_en = R0_en & R0_addr_sel == 8'hf7;
  assign mem_247_0_W0_addr = W0_addr[25:0];
  assign mem_247_0_W0_clk = W0_clk;
  assign mem_247_0_W0_data = W0_data[7:0];
  assign mem_247_0_W0_en = W0_en & W0_addr_sel == 8'hf7;
  assign mem_247_0_W0_mask = W0_mask[0];
  assign mem_247_1_R0_addr = R0_addr[25:0];
  assign mem_247_1_R0_clk = R0_clk;
  assign mem_247_1_R0_en = R0_en & R0_addr_sel == 8'hf7;
  assign mem_247_1_W0_addr = W0_addr[25:0];
  assign mem_247_1_W0_clk = W0_clk;
  assign mem_247_1_W0_data = W0_data[15:8];
  assign mem_247_1_W0_en = W0_en & W0_addr_sel == 8'hf7;
  assign mem_247_1_W0_mask = W0_mask[1];
  assign mem_247_2_R0_addr = R0_addr[25:0];
  assign mem_247_2_R0_clk = R0_clk;
  assign mem_247_2_R0_en = R0_en & R0_addr_sel == 8'hf7;
  assign mem_247_2_W0_addr = W0_addr[25:0];
  assign mem_247_2_W0_clk = W0_clk;
  assign mem_247_2_W0_data = W0_data[23:16];
  assign mem_247_2_W0_en = W0_en & W0_addr_sel == 8'hf7;
  assign mem_247_2_W0_mask = W0_mask[2];
  assign mem_247_3_R0_addr = R0_addr[25:0];
  assign mem_247_3_R0_clk = R0_clk;
  assign mem_247_3_R0_en = R0_en & R0_addr_sel == 8'hf7;
  assign mem_247_3_W0_addr = W0_addr[25:0];
  assign mem_247_3_W0_clk = W0_clk;
  assign mem_247_3_W0_data = W0_data[31:24];
  assign mem_247_3_W0_en = W0_en & W0_addr_sel == 8'hf7;
  assign mem_247_3_W0_mask = W0_mask[3];
  assign mem_247_4_R0_addr = R0_addr[25:0];
  assign mem_247_4_R0_clk = R0_clk;
  assign mem_247_4_R0_en = R0_en & R0_addr_sel == 8'hf7;
  assign mem_247_4_W0_addr = W0_addr[25:0];
  assign mem_247_4_W0_clk = W0_clk;
  assign mem_247_4_W0_data = W0_data[39:32];
  assign mem_247_4_W0_en = W0_en & W0_addr_sel == 8'hf7;
  assign mem_247_4_W0_mask = W0_mask[4];
  assign mem_247_5_R0_addr = R0_addr[25:0];
  assign mem_247_5_R0_clk = R0_clk;
  assign mem_247_5_R0_en = R0_en & R0_addr_sel == 8'hf7;
  assign mem_247_5_W0_addr = W0_addr[25:0];
  assign mem_247_5_W0_clk = W0_clk;
  assign mem_247_5_W0_data = W0_data[47:40];
  assign mem_247_5_W0_en = W0_en & W0_addr_sel == 8'hf7;
  assign mem_247_5_W0_mask = W0_mask[5];
  assign mem_247_6_R0_addr = R0_addr[25:0];
  assign mem_247_6_R0_clk = R0_clk;
  assign mem_247_6_R0_en = R0_en & R0_addr_sel == 8'hf7;
  assign mem_247_6_W0_addr = W0_addr[25:0];
  assign mem_247_6_W0_clk = W0_clk;
  assign mem_247_6_W0_data = W0_data[55:48];
  assign mem_247_6_W0_en = W0_en & W0_addr_sel == 8'hf7;
  assign mem_247_6_W0_mask = W0_mask[6];
  assign mem_247_7_R0_addr = R0_addr[25:0];
  assign mem_247_7_R0_clk = R0_clk;
  assign mem_247_7_R0_en = R0_en & R0_addr_sel == 8'hf7;
  assign mem_247_7_W0_addr = W0_addr[25:0];
  assign mem_247_7_W0_clk = W0_clk;
  assign mem_247_7_W0_data = W0_data[63:56];
  assign mem_247_7_W0_en = W0_en & W0_addr_sel == 8'hf7;
  assign mem_247_7_W0_mask = W0_mask[7];
  assign mem_248_0_R0_addr = R0_addr[25:0];
  assign mem_248_0_R0_clk = R0_clk;
  assign mem_248_0_R0_en = R0_en & R0_addr_sel == 8'hf8;
  assign mem_248_0_W0_addr = W0_addr[25:0];
  assign mem_248_0_W0_clk = W0_clk;
  assign mem_248_0_W0_data = W0_data[7:0];
  assign mem_248_0_W0_en = W0_en & W0_addr_sel == 8'hf8;
  assign mem_248_0_W0_mask = W0_mask[0];
  assign mem_248_1_R0_addr = R0_addr[25:0];
  assign mem_248_1_R0_clk = R0_clk;
  assign mem_248_1_R0_en = R0_en & R0_addr_sel == 8'hf8;
  assign mem_248_1_W0_addr = W0_addr[25:0];
  assign mem_248_1_W0_clk = W0_clk;
  assign mem_248_1_W0_data = W0_data[15:8];
  assign mem_248_1_W0_en = W0_en & W0_addr_sel == 8'hf8;
  assign mem_248_1_W0_mask = W0_mask[1];
  assign mem_248_2_R0_addr = R0_addr[25:0];
  assign mem_248_2_R0_clk = R0_clk;
  assign mem_248_2_R0_en = R0_en & R0_addr_sel == 8'hf8;
  assign mem_248_2_W0_addr = W0_addr[25:0];
  assign mem_248_2_W0_clk = W0_clk;
  assign mem_248_2_W0_data = W0_data[23:16];
  assign mem_248_2_W0_en = W0_en & W0_addr_sel == 8'hf8;
  assign mem_248_2_W0_mask = W0_mask[2];
  assign mem_248_3_R0_addr = R0_addr[25:0];
  assign mem_248_3_R0_clk = R0_clk;
  assign mem_248_3_R0_en = R0_en & R0_addr_sel == 8'hf8;
  assign mem_248_3_W0_addr = W0_addr[25:0];
  assign mem_248_3_W0_clk = W0_clk;
  assign mem_248_3_W0_data = W0_data[31:24];
  assign mem_248_3_W0_en = W0_en & W0_addr_sel == 8'hf8;
  assign mem_248_3_W0_mask = W0_mask[3];
  assign mem_248_4_R0_addr = R0_addr[25:0];
  assign mem_248_4_R0_clk = R0_clk;
  assign mem_248_4_R0_en = R0_en & R0_addr_sel == 8'hf8;
  assign mem_248_4_W0_addr = W0_addr[25:0];
  assign mem_248_4_W0_clk = W0_clk;
  assign mem_248_4_W0_data = W0_data[39:32];
  assign mem_248_4_W0_en = W0_en & W0_addr_sel == 8'hf8;
  assign mem_248_4_W0_mask = W0_mask[4];
  assign mem_248_5_R0_addr = R0_addr[25:0];
  assign mem_248_5_R0_clk = R0_clk;
  assign mem_248_5_R0_en = R0_en & R0_addr_sel == 8'hf8;
  assign mem_248_5_W0_addr = W0_addr[25:0];
  assign mem_248_5_W0_clk = W0_clk;
  assign mem_248_5_W0_data = W0_data[47:40];
  assign mem_248_5_W0_en = W0_en & W0_addr_sel == 8'hf8;
  assign mem_248_5_W0_mask = W0_mask[5];
  assign mem_248_6_R0_addr = R0_addr[25:0];
  assign mem_248_6_R0_clk = R0_clk;
  assign mem_248_6_R0_en = R0_en & R0_addr_sel == 8'hf8;
  assign mem_248_6_W0_addr = W0_addr[25:0];
  assign mem_248_6_W0_clk = W0_clk;
  assign mem_248_6_W0_data = W0_data[55:48];
  assign mem_248_6_W0_en = W0_en & W0_addr_sel == 8'hf8;
  assign mem_248_6_W0_mask = W0_mask[6];
  assign mem_248_7_R0_addr = R0_addr[25:0];
  assign mem_248_7_R0_clk = R0_clk;
  assign mem_248_7_R0_en = R0_en & R0_addr_sel == 8'hf8;
  assign mem_248_7_W0_addr = W0_addr[25:0];
  assign mem_248_7_W0_clk = W0_clk;
  assign mem_248_7_W0_data = W0_data[63:56];
  assign mem_248_7_W0_en = W0_en & W0_addr_sel == 8'hf8;
  assign mem_248_7_W0_mask = W0_mask[7];
  assign mem_249_0_R0_addr = R0_addr[25:0];
  assign mem_249_0_R0_clk = R0_clk;
  assign mem_249_0_R0_en = R0_en & R0_addr_sel == 8'hf9;
  assign mem_249_0_W0_addr = W0_addr[25:0];
  assign mem_249_0_W0_clk = W0_clk;
  assign mem_249_0_W0_data = W0_data[7:0];
  assign mem_249_0_W0_en = W0_en & W0_addr_sel == 8'hf9;
  assign mem_249_0_W0_mask = W0_mask[0];
  assign mem_249_1_R0_addr = R0_addr[25:0];
  assign mem_249_1_R0_clk = R0_clk;
  assign mem_249_1_R0_en = R0_en & R0_addr_sel == 8'hf9;
  assign mem_249_1_W0_addr = W0_addr[25:0];
  assign mem_249_1_W0_clk = W0_clk;
  assign mem_249_1_W0_data = W0_data[15:8];
  assign mem_249_1_W0_en = W0_en & W0_addr_sel == 8'hf9;
  assign mem_249_1_W0_mask = W0_mask[1];
  assign mem_249_2_R0_addr = R0_addr[25:0];
  assign mem_249_2_R0_clk = R0_clk;
  assign mem_249_2_R0_en = R0_en & R0_addr_sel == 8'hf9;
  assign mem_249_2_W0_addr = W0_addr[25:0];
  assign mem_249_2_W0_clk = W0_clk;
  assign mem_249_2_W0_data = W0_data[23:16];
  assign mem_249_2_W0_en = W0_en & W0_addr_sel == 8'hf9;
  assign mem_249_2_W0_mask = W0_mask[2];
  assign mem_249_3_R0_addr = R0_addr[25:0];
  assign mem_249_3_R0_clk = R0_clk;
  assign mem_249_3_R0_en = R0_en & R0_addr_sel == 8'hf9;
  assign mem_249_3_W0_addr = W0_addr[25:0];
  assign mem_249_3_W0_clk = W0_clk;
  assign mem_249_3_W0_data = W0_data[31:24];
  assign mem_249_3_W0_en = W0_en & W0_addr_sel == 8'hf9;
  assign mem_249_3_W0_mask = W0_mask[3];
  assign mem_249_4_R0_addr = R0_addr[25:0];
  assign mem_249_4_R0_clk = R0_clk;
  assign mem_249_4_R0_en = R0_en & R0_addr_sel == 8'hf9;
  assign mem_249_4_W0_addr = W0_addr[25:0];
  assign mem_249_4_W0_clk = W0_clk;
  assign mem_249_4_W0_data = W0_data[39:32];
  assign mem_249_4_W0_en = W0_en & W0_addr_sel == 8'hf9;
  assign mem_249_4_W0_mask = W0_mask[4];
  assign mem_249_5_R0_addr = R0_addr[25:0];
  assign mem_249_5_R0_clk = R0_clk;
  assign mem_249_5_R0_en = R0_en & R0_addr_sel == 8'hf9;
  assign mem_249_5_W0_addr = W0_addr[25:0];
  assign mem_249_5_W0_clk = W0_clk;
  assign mem_249_5_W0_data = W0_data[47:40];
  assign mem_249_5_W0_en = W0_en & W0_addr_sel == 8'hf9;
  assign mem_249_5_W0_mask = W0_mask[5];
  assign mem_249_6_R0_addr = R0_addr[25:0];
  assign mem_249_6_R0_clk = R0_clk;
  assign mem_249_6_R0_en = R0_en & R0_addr_sel == 8'hf9;
  assign mem_249_6_W0_addr = W0_addr[25:0];
  assign mem_249_6_W0_clk = W0_clk;
  assign mem_249_6_W0_data = W0_data[55:48];
  assign mem_249_6_W0_en = W0_en & W0_addr_sel == 8'hf9;
  assign mem_249_6_W0_mask = W0_mask[6];
  assign mem_249_7_R0_addr = R0_addr[25:0];
  assign mem_249_7_R0_clk = R0_clk;
  assign mem_249_7_R0_en = R0_en & R0_addr_sel == 8'hf9;
  assign mem_249_7_W0_addr = W0_addr[25:0];
  assign mem_249_7_W0_clk = W0_clk;
  assign mem_249_7_W0_data = W0_data[63:56];
  assign mem_249_7_W0_en = W0_en & W0_addr_sel == 8'hf9;
  assign mem_249_7_W0_mask = W0_mask[7];
  assign mem_250_0_R0_addr = R0_addr[25:0];
  assign mem_250_0_R0_clk = R0_clk;
  assign mem_250_0_R0_en = R0_en & R0_addr_sel == 8'hfa;
  assign mem_250_0_W0_addr = W0_addr[25:0];
  assign mem_250_0_W0_clk = W0_clk;
  assign mem_250_0_W0_data = W0_data[7:0];
  assign mem_250_0_W0_en = W0_en & W0_addr_sel == 8'hfa;
  assign mem_250_0_W0_mask = W0_mask[0];
  assign mem_250_1_R0_addr = R0_addr[25:0];
  assign mem_250_1_R0_clk = R0_clk;
  assign mem_250_1_R0_en = R0_en & R0_addr_sel == 8'hfa;
  assign mem_250_1_W0_addr = W0_addr[25:0];
  assign mem_250_1_W0_clk = W0_clk;
  assign mem_250_1_W0_data = W0_data[15:8];
  assign mem_250_1_W0_en = W0_en & W0_addr_sel == 8'hfa;
  assign mem_250_1_W0_mask = W0_mask[1];
  assign mem_250_2_R0_addr = R0_addr[25:0];
  assign mem_250_2_R0_clk = R0_clk;
  assign mem_250_2_R0_en = R0_en & R0_addr_sel == 8'hfa;
  assign mem_250_2_W0_addr = W0_addr[25:0];
  assign mem_250_2_W0_clk = W0_clk;
  assign mem_250_2_W0_data = W0_data[23:16];
  assign mem_250_2_W0_en = W0_en & W0_addr_sel == 8'hfa;
  assign mem_250_2_W0_mask = W0_mask[2];
  assign mem_250_3_R0_addr = R0_addr[25:0];
  assign mem_250_3_R0_clk = R0_clk;
  assign mem_250_3_R0_en = R0_en & R0_addr_sel == 8'hfa;
  assign mem_250_3_W0_addr = W0_addr[25:0];
  assign mem_250_3_W0_clk = W0_clk;
  assign mem_250_3_W0_data = W0_data[31:24];
  assign mem_250_3_W0_en = W0_en & W0_addr_sel == 8'hfa;
  assign mem_250_3_W0_mask = W0_mask[3];
  assign mem_250_4_R0_addr = R0_addr[25:0];
  assign mem_250_4_R0_clk = R0_clk;
  assign mem_250_4_R0_en = R0_en & R0_addr_sel == 8'hfa;
  assign mem_250_4_W0_addr = W0_addr[25:0];
  assign mem_250_4_W0_clk = W0_clk;
  assign mem_250_4_W0_data = W0_data[39:32];
  assign mem_250_4_W0_en = W0_en & W0_addr_sel == 8'hfa;
  assign mem_250_4_W0_mask = W0_mask[4];
  assign mem_250_5_R0_addr = R0_addr[25:0];
  assign mem_250_5_R0_clk = R0_clk;
  assign mem_250_5_R0_en = R0_en & R0_addr_sel == 8'hfa;
  assign mem_250_5_W0_addr = W0_addr[25:0];
  assign mem_250_5_W0_clk = W0_clk;
  assign mem_250_5_W0_data = W0_data[47:40];
  assign mem_250_5_W0_en = W0_en & W0_addr_sel == 8'hfa;
  assign mem_250_5_W0_mask = W0_mask[5];
  assign mem_250_6_R0_addr = R0_addr[25:0];
  assign mem_250_6_R0_clk = R0_clk;
  assign mem_250_6_R0_en = R0_en & R0_addr_sel == 8'hfa;
  assign mem_250_6_W0_addr = W0_addr[25:0];
  assign mem_250_6_W0_clk = W0_clk;
  assign mem_250_6_W0_data = W0_data[55:48];
  assign mem_250_6_W0_en = W0_en & W0_addr_sel == 8'hfa;
  assign mem_250_6_W0_mask = W0_mask[6];
  assign mem_250_7_R0_addr = R0_addr[25:0];
  assign mem_250_7_R0_clk = R0_clk;
  assign mem_250_7_R0_en = R0_en & R0_addr_sel == 8'hfa;
  assign mem_250_7_W0_addr = W0_addr[25:0];
  assign mem_250_7_W0_clk = W0_clk;
  assign mem_250_7_W0_data = W0_data[63:56];
  assign mem_250_7_W0_en = W0_en & W0_addr_sel == 8'hfa;
  assign mem_250_7_W0_mask = W0_mask[7];
  assign mem_251_0_R0_addr = R0_addr[25:0];
  assign mem_251_0_R0_clk = R0_clk;
  assign mem_251_0_R0_en = R0_en & R0_addr_sel == 8'hfb;
  assign mem_251_0_W0_addr = W0_addr[25:0];
  assign mem_251_0_W0_clk = W0_clk;
  assign mem_251_0_W0_data = W0_data[7:0];
  assign mem_251_0_W0_en = W0_en & W0_addr_sel == 8'hfb;
  assign mem_251_0_W0_mask = W0_mask[0];
  assign mem_251_1_R0_addr = R0_addr[25:0];
  assign mem_251_1_R0_clk = R0_clk;
  assign mem_251_1_R0_en = R0_en & R0_addr_sel == 8'hfb;
  assign mem_251_1_W0_addr = W0_addr[25:0];
  assign mem_251_1_W0_clk = W0_clk;
  assign mem_251_1_W0_data = W0_data[15:8];
  assign mem_251_1_W0_en = W0_en & W0_addr_sel == 8'hfb;
  assign mem_251_1_W0_mask = W0_mask[1];
  assign mem_251_2_R0_addr = R0_addr[25:0];
  assign mem_251_2_R0_clk = R0_clk;
  assign mem_251_2_R0_en = R0_en & R0_addr_sel == 8'hfb;
  assign mem_251_2_W0_addr = W0_addr[25:0];
  assign mem_251_2_W0_clk = W0_clk;
  assign mem_251_2_W0_data = W0_data[23:16];
  assign mem_251_2_W0_en = W0_en & W0_addr_sel == 8'hfb;
  assign mem_251_2_W0_mask = W0_mask[2];
  assign mem_251_3_R0_addr = R0_addr[25:0];
  assign mem_251_3_R0_clk = R0_clk;
  assign mem_251_3_R0_en = R0_en & R0_addr_sel == 8'hfb;
  assign mem_251_3_W0_addr = W0_addr[25:0];
  assign mem_251_3_W0_clk = W0_clk;
  assign mem_251_3_W0_data = W0_data[31:24];
  assign mem_251_3_W0_en = W0_en & W0_addr_sel == 8'hfb;
  assign mem_251_3_W0_mask = W0_mask[3];
  assign mem_251_4_R0_addr = R0_addr[25:0];
  assign mem_251_4_R0_clk = R0_clk;
  assign mem_251_4_R0_en = R0_en & R0_addr_sel == 8'hfb;
  assign mem_251_4_W0_addr = W0_addr[25:0];
  assign mem_251_4_W0_clk = W0_clk;
  assign mem_251_4_W0_data = W0_data[39:32];
  assign mem_251_4_W0_en = W0_en & W0_addr_sel == 8'hfb;
  assign mem_251_4_W0_mask = W0_mask[4];
  assign mem_251_5_R0_addr = R0_addr[25:0];
  assign mem_251_5_R0_clk = R0_clk;
  assign mem_251_5_R0_en = R0_en & R0_addr_sel == 8'hfb;
  assign mem_251_5_W0_addr = W0_addr[25:0];
  assign mem_251_5_W0_clk = W0_clk;
  assign mem_251_5_W0_data = W0_data[47:40];
  assign mem_251_5_W0_en = W0_en & W0_addr_sel == 8'hfb;
  assign mem_251_5_W0_mask = W0_mask[5];
  assign mem_251_6_R0_addr = R0_addr[25:0];
  assign mem_251_6_R0_clk = R0_clk;
  assign mem_251_6_R0_en = R0_en & R0_addr_sel == 8'hfb;
  assign mem_251_6_W0_addr = W0_addr[25:0];
  assign mem_251_6_W0_clk = W0_clk;
  assign mem_251_6_W0_data = W0_data[55:48];
  assign mem_251_6_W0_en = W0_en & W0_addr_sel == 8'hfb;
  assign mem_251_6_W0_mask = W0_mask[6];
  assign mem_251_7_R0_addr = R0_addr[25:0];
  assign mem_251_7_R0_clk = R0_clk;
  assign mem_251_7_R0_en = R0_en & R0_addr_sel == 8'hfb;
  assign mem_251_7_W0_addr = W0_addr[25:0];
  assign mem_251_7_W0_clk = W0_clk;
  assign mem_251_7_W0_data = W0_data[63:56];
  assign mem_251_7_W0_en = W0_en & W0_addr_sel == 8'hfb;
  assign mem_251_7_W0_mask = W0_mask[7];
  assign mem_252_0_R0_addr = R0_addr[25:0];
  assign mem_252_0_R0_clk = R0_clk;
  assign mem_252_0_R0_en = R0_en & R0_addr_sel == 8'hfc;
  assign mem_252_0_W0_addr = W0_addr[25:0];
  assign mem_252_0_W0_clk = W0_clk;
  assign mem_252_0_W0_data = W0_data[7:0];
  assign mem_252_0_W0_en = W0_en & W0_addr_sel == 8'hfc;
  assign mem_252_0_W0_mask = W0_mask[0];
  assign mem_252_1_R0_addr = R0_addr[25:0];
  assign mem_252_1_R0_clk = R0_clk;
  assign mem_252_1_R0_en = R0_en & R0_addr_sel == 8'hfc;
  assign mem_252_1_W0_addr = W0_addr[25:0];
  assign mem_252_1_W0_clk = W0_clk;
  assign mem_252_1_W0_data = W0_data[15:8];
  assign mem_252_1_W0_en = W0_en & W0_addr_sel == 8'hfc;
  assign mem_252_1_W0_mask = W0_mask[1];
  assign mem_252_2_R0_addr = R0_addr[25:0];
  assign mem_252_2_R0_clk = R0_clk;
  assign mem_252_2_R0_en = R0_en & R0_addr_sel == 8'hfc;
  assign mem_252_2_W0_addr = W0_addr[25:0];
  assign mem_252_2_W0_clk = W0_clk;
  assign mem_252_2_W0_data = W0_data[23:16];
  assign mem_252_2_W0_en = W0_en & W0_addr_sel == 8'hfc;
  assign mem_252_2_W0_mask = W0_mask[2];
  assign mem_252_3_R0_addr = R0_addr[25:0];
  assign mem_252_3_R0_clk = R0_clk;
  assign mem_252_3_R0_en = R0_en & R0_addr_sel == 8'hfc;
  assign mem_252_3_W0_addr = W0_addr[25:0];
  assign mem_252_3_W0_clk = W0_clk;
  assign mem_252_3_W0_data = W0_data[31:24];
  assign mem_252_3_W0_en = W0_en & W0_addr_sel == 8'hfc;
  assign mem_252_3_W0_mask = W0_mask[3];
  assign mem_252_4_R0_addr = R0_addr[25:0];
  assign mem_252_4_R0_clk = R0_clk;
  assign mem_252_4_R0_en = R0_en & R0_addr_sel == 8'hfc;
  assign mem_252_4_W0_addr = W0_addr[25:0];
  assign mem_252_4_W0_clk = W0_clk;
  assign mem_252_4_W0_data = W0_data[39:32];
  assign mem_252_4_W0_en = W0_en & W0_addr_sel == 8'hfc;
  assign mem_252_4_W0_mask = W0_mask[4];
  assign mem_252_5_R0_addr = R0_addr[25:0];
  assign mem_252_5_R0_clk = R0_clk;
  assign mem_252_5_R0_en = R0_en & R0_addr_sel == 8'hfc;
  assign mem_252_5_W0_addr = W0_addr[25:0];
  assign mem_252_5_W0_clk = W0_clk;
  assign mem_252_5_W0_data = W0_data[47:40];
  assign mem_252_5_W0_en = W0_en & W0_addr_sel == 8'hfc;
  assign mem_252_5_W0_mask = W0_mask[5];
  assign mem_252_6_R0_addr = R0_addr[25:0];
  assign mem_252_6_R0_clk = R0_clk;
  assign mem_252_6_R0_en = R0_en & R0_addr_sel == 8'hfc;
  assign mem_252_6_W0_addr = W0_addr[25:0];
  assign mem_252_6_W0_clk = W0_clk;
  assign mem_252_6_W0_data = W0_data[55:48];
  assign mem_252_6_W0_en = W0_en & W0_addr_sel == 8'hfc;
  assign mem_252_6_W0_mask = W0_mask[6];
  assign mem_252_7_R0_addr = R0_addr[25:0];
  assign mem_252_7_R0_clk = R0_clk;
  assign mem_252_7_R0_en = R0_en & R0_addr_sel == 8'hfc;
  assign mem_252_7_W0_addr = W0_addr[25:0];
  assign mem_252_7_W0_clk = W0_clk;
  assign mem_252_7_W0_data = W0_data[63:56];
  assign mem_252_7_W0_en = W0_en & W0_addr_sel == 8'hfc;
  assign mem_252_7_W0_mask = W0_mask[7];
  assign mem_253_0_R0_addr = R0_addr[25:0];
  assign mem_253_0_R0_clk = R0_clk;
  assign mem_253_0_R0_en = R0_en & R0_addr_sel == 8'hfd;
  assign mem_253_0_W0_addr = W0_addr[25:0];
  assign mem_253_0_W0_clk = W0_clk;
  assign mem_253_0_W0_data = W0_data[7:0];
  assign mem_253_0_W0_en = W0_en & W0_addr_sel == 8'hfd;
  assign mem_253_0_W0_mask = W0_mask[0];
  assign mem_253_1_R0_addr = R0_addr[25:0];
  assign mem_253_1_R0_clk = R0_clk;
  assign mem_253_1_R0_en = R0_en & R0_addr_sel == 8'hfd;
  assign mem_253_1_W0_addr = W0_addr[25:0];
  assign mem_253_1_W0_clk = W0_clk;
  assign mem_253_1_W0_data = W0_data[15:8];
  assign mem_253_1_W0_en = W0_en & W0_addr_sel == 8'hfd;
  assign mem_253_1_W0_mask = W0_mask[1];
  assign mem_253_2_R0_addr = R0_addr[25:0];
  assign mem_253_2_R0_clk = R0_clk;
  assign mem_253_2_R0_en = R0_en & R0_addr_sel == 8'hfd;
  assign mem_253_2_W0_addr = W0_addr[25:0];
  assign mem_253_2_W0_clk = W0_clk;
  assign mem_253_2_W0_data = W0_data[23:16];
  assign mem_253_2_W0_en = W0_en & W0_addr_sel == 8'hfd;
  assign mem_253_2_W0_mask = W0_mask[2];
  assign mem_253_3_R0_addr = R0_addr[25:0];
  assign mem_253_3_R0_clk = R0_clk;
  assign mem_253_3_R0_en = R0_en & R0_addr_sel == 8'hfd;
  assign mem_253_3_W0_addr = W0_addr[25:0];
  assign mem_253_3_W0_clk = W0_clk;
  assign mem_253_3_W0_data = W0_data[31:24];
  assign mem_253_3_W0_en = W0_en & W0_addr_sel == 8'hfd;
  assign mem_253_3_W0_mask = W0_mask[3];
  assign mem_253_4_R0_addr = R0_addr[25:0];
  assign mem_253_4_R0_clk = R0_clk;
  assign mem_253_4_R0_en = R0_en & R0_addr_sel == 8'hfd;
  assign mem_253_4_W0_addr = W0_addr[25:0];
  assign mem_253_4_W0_clk = W0_clk;
  assign mem_253_4_W0_data = W0_data[39:32];
  assign mem_253_4_W0_en = W0_en & W0_addr_sel == 8'hfd;
  assign mem_253_4_W0_mask = W0_mask[4];
  assign mem_253_5_R0_addr = R0_addr[25:0];
  assign mem_253_5_R0_clk = R0_clk;
  assign mem_253_5_R0_en = R0_en & R0_addr_sel == 8'hfd;
  assign mem_253_5_W0_addr = W0_addr[25:0];
  assign mem_253_5_W0_clk = W0_clk;
  assign mem_253_5_W0_data = W0_data[47:40];
  assign mem_253_5_W0_en = W0_en & W0_addr_sel == 8'hfd;
  assign mem_253_5_W0_mask = W0_mask[5];
  assign mem_253_6_R0_addr = R0_addr[25:0];
  assign mem_253_6_R0_clk = R0_clk;
  assign mem_253_6_R0_en = R0_en & R0_addr_sel == 8'hfd;
  assign mem_253_6_W0_addr = W0_addr[25:0];
  assign mem_253_6_W0_clk = W0_clk;
  assign mem_253_6_W0_data = W0_data[55:48];
  assign mem_253_6_W0_en = W0_en & W0_addr_sel == 8'hfd;
  assign mem_253_6_W0_mask = W0_mask[6];
  assign mem_253_7_R0_addr = R0_addr[25:0];
  assign mem_253_7_R0_clk = R0_clk;
  assign mem_253_7_R0_en = R0_en & R0_addr_sel == 8'hfd;
  assign mem_253_7_W0_addr = W0_addr[25:0];
  assign mem_253_7_W0_clk = W0_clk;
  assign mem_253_7_W0_data = W0_data[63:56];
  assign mem_253_7_W0_en = W0_en & W0_addr_sel == 8'hfd;
  assign mem_253_7_W0_mask = W0_mask[7];
  assign mem_254_0_R0_addr = R0_addr[25:0];
  assign mem_254_0_R0_clk = R0_clk;
  assign mem_254_0_R0_en = R0_en & R0_addr_sel == 8'hfe;
  assign mem_254_0_W0_addr = W0_addr[25:0];
  assign mem_254_0_W0_clk = W0_clk;
  assign mem_254_0_W0_data = W0_data[7:0];
  assign mem_254_0_W0_en = W0_en & W0_addr_sel == 8'hfe;
  assign mem_254_0_W0_mask = W0_mask[0];
  assign mem_254_1_R0_addr = R0_addr[25:0];
  assign mem_254_1_R0_clk = R0_clk;
  assign mem_254_1_R0_en = R0_en & R0_addr_sel == 8'hfe;
  assign mem_254_1_W0_addr = W0_addr[25:0];
  assign mem_254_1_W0_clk = W0_clk;
  assign mem_254_1_W0_data = W0_data[15:8];
  assign mem_254_1_W0_en = W0_en & W0_addr_sel == 8'hfe;
  assign mem_254_1_W0_mask = W0_mask[1];
  assign mem_254_2_R0_addr = R0_addr[25:0];
  assign mem_254_2_R0_clk = R0_clk;
  assign mem_254_2_R0_en = R0_en & R0_addr_sel == 8'hfe;
  assign mem_254_2_W0_addr = W0_addr[25:0];
  assign mem_254_2_W0_clk = W0_clk;
  assign mem_254_2_W0_data = W0_data[23:16];
  assign mem_254_2_W0_en = W0_en & W0_addr_sel == 8'hfe;
  assign mem_254_2_W0_mask = W0_mask[2];
  assign mem_254_3_R0_addr = R0_addr[25:0];
  assign mem_254_3_R0_clk = R0_clk;
  assign mem_254_3_R0_en = R0_en & R0_addr_sel == 8'hfe;
  assign mem_254_3_W0_addr = W0_addr[25:0];
  assign mem_254_3_W0_clk = W0_clk;
  assign mem_254_3_W0_data = W0_data[31:24];
  assign mem_254_3_W0_en = W0_en & W0_addr_sel == 8'hfe;
  assign mem_254_3_W0_mask = W0_mask[3];
  assign mem_254_4_R0_addr = R0_addr[25:0];
  assign mem_254_4_R0_clk = R0_clk;
  assign mem_254_4_R0_en = R0_en & R0_addr_sel == 8'hfe;
  assign mem_254_4_W0_addr = W0_addr[25:0];
  assign mem_254_4_W0_clk = W0_clk;
  assign mem_254_4_W0_data = W0_data[39:32];
  assign mem_254_4_W0_en = W0_en & W0_addr_sel == 8'hfe;
  assign mem_254_4_W0_mask = W0_mask[4];
  assign mem_254_5_R0_addr = R0_addr[25:0];
  assign mem_254_5_R0_clk = R0_clk;
  assign mem_254_5_R0_en = R0_en & R0_addr_sel == 8'hfe;
  assign mem_254_5_W0_addr = W0_addr[25:0];
  assign mem_254_5_W0_clk = W0_clk;
  assign mem_254_5_W0_data = W0_data[47:40];
  assign mem_254_5_W0_en = W0_en & W0_addr_sel == 8'hfe;
  assign mem_254_5_W0_mask = W0_mask[5];
  assign mem_254_6_R0_addr = R0_addr[25:0];
  assign mem_254_6_R0_clk = R0_clk;
  assign mem_254_6_R0_en = R0_en & R0_addr_sel == 8'hfe;
  assign mem_254_6_W0_addr = W0_addr[25:0];
  assign mem_254_6_W0_clk = W0_clk;
  assign mem_254_6_W0_data = W0_data[55:48];
  assign mem_254_6_W0_en = W0_en & W0_addr_sel == 8'hfe;
  assign mem_254_6_W0_mask = W0_mask[6];
  assign mem_254_7_R0_addr = R0_addr[25:0];
  assign mem_254_7_R0_clk = R0_clk;
  assign mem_254_7_R0_en = R0_en & R0_addr_sel == 8'hfe;
  assign mem_254_7_W0_addr = W0_addr[25:0];
  assign mem_254_7_W0_clk = W0_clk;
  assign mem_254_7_W0_data = W0_data[63:56];
  assign mem_254_7_W0_en = W0_en & W0_addr_sel == 8'hfe;
  assign mem_254_7_W0_mask = W0_mask[7];
  assign mem_255_0_R0_addr = R0_addr[25:0];
  assign mem_255_0_R0_clk = R0_clk;
  assign mem_255_0_R0_en = R0_en & R0_addr_sel == 8'hff;
  assign mem_255_0_W0_addr = W0_addr[25:0];
  assign mem_255_0_W0_clk = W0_clk;
  assign mem_255_0_W0_data = W0_data[7:0];
  assign mem_255_0_W0_en = W0_en & W0_addr_sel == 8'hff;
  assign mem_255_0_W0_mask = W0_mask[0];
  assign mem_255_1_R0_addr = R0_addr[25:0];
  assign mem_255_1_R0_clk = R0_clk;
  assign mem_255_1_R0_en = R0_en & R0_addr_sel == 8'hff;
  assign mem_255_1_W0_addr = W0_addr[25:0];
  assign mem_255_1_W0_clk = W0_clk;
  assign mem_255_1_W0_data = W0_data[15:8];
  assign mem_255_1_W0_en = W0_en & W0_addr_sel == 8'hff;
  assign mem_255_1_W0_mask = W0_mask[1];
  assign mem_255_2_R0_addr = R0_addr[25:0];
  assign mem_255_2_R0_clk = R0_clk;
  assign mem_255_2_R0_en = R0_en & R0_addr_sel == 8'hff;
  assign mem_255_2_W0_addr = W0_addr[25:0];
  assign mem_255_2_W0_clk = W0_clk;
  assign mem_255_2_W0_data = W0_data[23:16];
  assign mem_255_2_W0_en = W0_en & W0_addr_sel == 8'hff;
  assign mem_255_2_W0_mask = W0_mask[2];
  assign mem_255_3_R0_addr = R0_addr[25:0];
  assign mem_255_3_R0_clk = R0_clk;
  assign mem_255_3_R0_en = R0_en & R0_addr_sel == 8'hff;
  assign mem_255_3_W0_addr = W0_addr[25:0];
  assign mem_255_3_W0_clk = W0_clk;
  assign mem_255_3_W0_data = W0_data[31:24];
  assign mem_255_3_W0_en = W0_en & W0_addr_sel == 8'hff;
  assign mem_255_3_W0_mask = W0_mask[3];
  assign mem_255_4_R0_addr = R0_addr[25:0];
  assign mem_255_4_R0_clk = R0_clk;
  assign mem_255_4_R0_en = R0_en & R0_addr_sel == 8'hff;
  assign mem_255_4_W0_addr = W0_addr[25:0];
  assign mem_255_4_W0_clk = W0_clk;
  assign mem_255_4_W0_data = W0_data[39:32];
  assign mem_255_4_W0_en = W0_en & W0_addr_sel == 8'hff;
  assign mem_255_4_W0_mask = W0_mask[4];
  assign mem_255_5_R0_addr = R0_addr[25:0];
  assign mem_255_5_R0_clk = R0_clk;
  assign mem_255_5_R0_en = R0_en & R0_addr_sel == 8'hff;
  assign mem_255_5_W0_addr = W0_addr[25:0];
  assign mem_255_5_W0_clk = W0_clk;
  assign mem_255_5_W0_data = W0_data[47:40];
  assign mem_255_5_W0_en = W0_en & W0_addr_sel == 8'hff;
  assign mem_255_5_W0_mask = W0_mask[5];
  assign mem_255_6_R0_addr = R0_addr[25:0];
  assign mem_255_6_R0_clk = R0_clk;
  assign mem_255_6_R0_en = R0_en & R0_addr_sel == 8'hff;
  assign mem_255_6_W0_addr = W0_addr[25:0];
  assign mem_255_6_W0_clk = W0_clk;
  assign mem_255_6_W0_data = W0_data[55:48];
  assign mem_255_6_W0_en = W0_en & W0_addr_sel == 8'hff;
  assign mem_255_6_W0_mask = W0_mask[6];
  assign mem_255_7_R0_addr = R0_addr[25:0];
  assign mem_255_7_R0_clk = R0_clk;
  assign mem_255_7_R0_en = R0_en & R0_addr_sel == 8'hff;
  assign mem_255_7_W0_addr = W0_addr[25:0];
  assign mem_255_7_W0_clk = W0_clk;
  assign mem_255_7_W0_data = W0_data[63:56];
  assign mem_255_7_W0_en = W0_en & W0_addr_sel == 8'hff;
  assign mem_255_7_W0_mask = W0_mask[7];
  always @(posedge R0_clk) begin
    if (R0_en) begin
      R0_addr_sel_reg <= R0_addr_sel;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  R0_addr_sel_reg = _RAND_0[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule

module split_mem_0_ext(
  input  [25:0] R0_addr,
  input         R0_clk,
  output [7:0]  R0_data,
  input         R0_en,
  input  [25:0] W0_addr,
  input         W0_clk,
  input  [7:0]  W0_data,
  input         W0_en,
  input         W0_mask
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] ram [0:67108863];
  wire  ram_R_0_en;
  wire [25:0] ram_R_0_addr;
  wire [7:0] ram_R_0_data;
  wire [7:0] ram_W_0_data;
  wire [25:0] ram_W_0_addr;
  wire  ram_W_0_mask;
  wire  ram_W_0_en;
  reg  ram_R_0_en_pipe_0;
  reg [25:0] ram_R_0_addr_pipe_0;
  assign ram_R_0_en = ram_R_0_en_pipe_0;
  assign ram_R_0_addr = ram_R_0_addr_pipe_0;
  assign ram_R_0_data = ram[ram_R_0_addr];
  assign ram_W_0_data = W0_data;
  assign ram_W_0_addr = W0_addr;
  assign ram_W_0_mask = W0_mask;
  assign ram_W_0_en = W0_en;
  assign R0_data = ram_R_0_data;
  always @(posedge W0_clk) begin
    if (ram_W_0_en & ram_W_0_mask) begin
      ram[ram_W_0_addr] <= ram_W_0_data;
    end
  end
  always @(posedge R0_clk) begin
    ram_R_0_en_pipe_0 <= R0_en;
    if (R0_en) begin
      ram_R_0_addr_pipe_0 <= R0_addr;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 67108864; initvar = initvar+1)
    ram[initvar] = _RAND_0[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  ram_R_0_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  ram_R_0_addr_pipe_0 = _RAND_2[25:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
